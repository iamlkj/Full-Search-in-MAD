
module MC2_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X2 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHX1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MC2_DW01_sub_5 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [7:1] carry;

  ADDFXL U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFHX2 U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFX2 U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XNOR2XL U1 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[4]), .Y(n4) );
  INVXL U3 ( .A(B[2]), .Y(n6) );
  INVXL U4 ( .A(B[5]), .Y(n3) );
  INVXL U5 ( .A(B[3]), .Y(n5) );
  INVXL U6 ( .A(B[1]), .Y(n7) );
  INVXL U7 ( .A(A[0]), .Y(n1) );
  INVXL U8 ( .A(B[0]), .Y(n8) );
  INVXL U9 ( .A(B[6]), .Y(n2) );
  XNOR3XL U10 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(DIFF[7]) );
  NAND2X1 U11 ( .A(B[0]), .B(n1), .Y(carry[1]) );
endmodule


module MC2_DW01_sub_6 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [7:1] carry;

  ADDFXL U2_3 ( .A(A[3]), .B(n7), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n5), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  XOR3X1 U2_7 ( .A(A[7]), .B(n3), .C(carry[7]), .Y(DIFF[7]) );
  ADDFX2 U2_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n6), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFHX2 U2_1 ( .A(A[1]), .B(n9), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  ADDFHX1 U2_2 ( .A(A[2]), .B(n8), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  INVXL U1 ( .A(A[0]), .Y(n2) );
  XNOR2XL U2 ( .A(n10), .B(A[0]), .Y(DIFF[0]) );
  INVXL U3 ( .A(B[5]), .Y(n5) );
  INVXL U4 ( .A(B[3]), .Y(n7) );
  INVXL U5 ( .A(B[4]), .Y(n6) );
  INVXL U6 ( .A(B[2]), .Y(n8) );
  INVXL U7 ( .A(B[0]), .Y(n10) );
  INVXL U8 ( .A(B[6]), .Y(n4) );
  INVXL U9 ( .A(B[7]), .Y(n3) );
  CLKINVX1 U10 ( .A(n10), .Y(n1) );
  CLKINVX1 U11 ( .A(B[1]), .Y(n9) );
  NAND2X1 U12 ( .A(n1), .B(n2), .Y(carry[1]) );
endmodule


module MC2_DW01_sub_7 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [7:1] carry;

  ADDFXL U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XNOR3X1 U1 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(DIFF[7]) );
  INVXL U2 ( .A(B[0]), .Y(n8) );
  XNOR2XL U3 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVXL U4 ( .A(B[2]), .Y(n6) );
  INVXL U5 ( .A(B[4]), .Y(n4) );
  INVXL U6 ( .A(B[3]), .Y(n5) );
  INVXL U7 ( .A(B[1]), .Y(n7) );
  INVXL U8 ( .A(A[0]), .Y(n1) );
  INVXL U9 ( .A(B[6]), .Y(n2) );
  NAND2X1 U10 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U11 ( .A(B[5]), .Y(n3) );
endmodule


module MC2_DW01_sub_8 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  ADDFXL U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XOR3X1 U2_7 ( .A(A[7]), .B(n2), .C(carry[7]), .Y(DIFF[7]) );
  ADDFX2 U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XNOR2XL U1 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[3]), .Y(n6) );
  INVXL U3 ( .A(B[4]), .Y(n5) );
  INVXL U4 ( .A(B[2]), .Y(n7) );
  INVXL U5 ( .A(B[0]), .Y(n9) );
  INVXL U6 ( .A(B[6]), .Y(n3) );
  INVXL U7 ( .A(B[7]), .Y(n2) );
  CLKINVX1 U8 ( .A(B[5]), .Y(n4) );
  CLKINVX1 U9 ( .A(B[1]), .Y(n8) );
  NAND2X1 U10 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U11 ( .A(A[0]), .Y(n1) );
endmodule


module MC2_DW01_sub_9 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [7:1] carry;

  ADDFXL U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  XNOR2XL U1 ( .A(n8), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[4]), .Y(n4) );
  INVXL U3 ( .A(B[2]), .Y(n6) );
  INVXL U4 ( .A(B[5]), .Y(n3) );
  INVXL U5 ( .A(B[3]), .Y(n5) );
  INVXL U6 ( .A(B[1]), .Y(n7) );
  INVXL U7 ( .A(A[0]), .Y(n1) );
  INVXL U8 ( .A(B[0]), .Y(n8) );
  INVXL U9 ( .A(B[6]), .Y(n2) );
  XNOR3XL U10 ( .A(A[7]), .B(B[7]), .C(carry[7]), .Y(DIFF[7]) );
  NAND2X1 U11 ( .A(B[0]), .B(n1), .Y(carry[1]) );
endmodule


module MC2_DW01_sub_10 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  ADDFXL U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  XOR3X1 U2_7 ( .A(A[7]), .B(n2), .C(carry[7]), .Y(DIFF[7]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  ADDFX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  XNOR2XL U1 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[5]), .Y(n4) );
  INVXL U3 ( .A(B[3]), .Y(n6) );
  INVXL U4 ( .A(B[4]), .Y(n5) );
  INVXL U5 ( .A(B[2]), .Y(n7) );
  INVXL U6 ( .A(B[0]), .Y(n9) );
  INVXL U7 ( .A(B[6]), .Y(n3) );
  INVXL U8 ( .A(B[7]), .Y(n2) );
  CLKINVX1 U9 ( .A(B[1]), .Y(n8) );
  NAND2X1 U10 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U11 ( .A(A[0]), .Y(n1) );
endmodule


module MC2_DW01_sub_11 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  ADDFXL U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  ADDFXL U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XOR3X1 U2_7 ( .A(A[7]), .B(n2), .C(carry[7]), .Y(DIFF[7]) );
  XNOR2XL U1 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[7]), .Y(n2) );
  INVXL U3 ( .A(B[4]), .Y(n5) );
  INVXL U4 ( .A(B[2]), .Y(n7) );
  INVXL U5 ( .A(B[5]), .Y(n4) );
  INVXL U6 ( .A(B[3]), .Y(n6) );
  INVXL U7 ( .A(B[1]), .Y(n8) );
  INVXL U8 ( .A(A[0]), .Y(n1) );
  INVXL U9 ( .A(B[0]), .Y(n9) );
  INVXL U10 ( .A(B[6]), .Y(n3) );
  NAND2X1 U11 ( .A(B[0]), .B(n1), .Y(carry[1]) );
endmodule


module MC2_DW01_sub_12 ( A, B, DIFF );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:1] carry;

  ADDFXL U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  ADDFXL U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  ADDFXL U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  ADDFXL U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  XOR3X1 U2_7 ( .A(A[7]), .B(n2), .C(carry[7]), .Y(DIFF[7]) );
  ADDFHX2 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  ADDFX2 U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XNOR2XL U1 ( .A(n9), .B(A[0]), .Y(DIFF[0]) );
  INVXL U2 ( .A(B[5]), .Y(n4) );
  INVXL U3 ( .A(B[3]), .Y(n6) );
  INVXL U4 ( .A(B[4]), .Y(n5) );
  INVXL U5 ( .A(B[2]), .Y(n7) );
  INVXL U6 ( .A(B[0]), .Y(n9) );
  INVXL U7 ( .A(B[6]), .Y(n3) );
  INVXL U8 ( .A(B[7]), .Y(n2) );
  CLKINVX1 U9 ( .A(B[1]), .Y(n8) );
  NAND2X1 U10 ( .A(B[0]), .B(n1), .Y(carry[1]) );
  CLKINVX1 U11 ( .A(A[0]), .Y(n1) );
endmodule


module MC2_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MC2_DW01_add_5 ( A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, B_6_, B_5_, B_4_,
         B_3_, B_2_, B_1_, B_0_;
  output SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_,
         SUM_0_;
  wire   n1;
  wire   [7:2] carry;

  CMPR32X2 U1_7 ( .A(A_7_), .B(B_7_), .C(carry[7]), .CO(SUM_8_), .S(SUM_7_) );
  CMPR32X2 U1_6 ( .A(A_6_), .B(B_6_), .C(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  CMPR32X2 U1_5 ( .A(A_5_), .B(B_5_), .C(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFX1 U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  CMPR32X2 U1_4 ( .A(A_4_), .B(B_4_), .C(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFHX2 U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFX2 U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_add_4 ( A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, B_6_, B_5_, B_4_,
         B_3_, B_2_, B_1_, B_0_;
  output SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_,
         SUM_0_;
  wire   n1, n2, n3, n4;
  wire   [7:2] carry;

  ADDFHX1 U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFX1 U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  CMPR32X2 U1_4 ( .A(A_4_), .B(B_4_), .C(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFX1 U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFHX2 U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFX2 U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR3X1 U2 ( .A(carry[7]), .B(A_7_), .C(B_7_), .Y(SUM_7_) );
  NAND2X1 U3 ( .A(B_7_), .B(carry[7]), .Y(n2) );
  NAND2X1 U4 ( .A(A_7_), .B(carry[7]), .Y(n3) );
  NAND2X1 U5 ( .A(A_7_), .B(B_7_), .Y(n4) );
  NAND3X1 U6 ( .A(n2), .B(n3), .C(n4), .Y(SUM_8_) );
  XOR2X1 U7 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_add_3 ( A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, 
        B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_9_, SUM_8_, 
        SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_8_, B_7_, B_6_,
         B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_,
         SUM_1_, SUM_0_;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n1;

  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  ADDFHX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  CMPR32X2 U1_3 ( .A(A_3_), .B(B_3_), .C(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  ADDFX1 U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFHX2 U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  ADDFHX2 U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(SUM_9_), .S(SUM_8_) );
  ADDFX2 U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2XL U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_add_2 ( A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, B_6_, B_5_, B_4_,
         B_3_, B_2_, B_1_, B_0_;
  output SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_,
         SUM_0_;
  wire   n1;
  wire   [7:2] carry;

  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(SUM_8_), .S(SUM_7_) );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_add_1 ( A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, 
        B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_7_, B_6_, B_5_, B_4_,
         B_3_, B_2_, B_1_, B_0_;
  output SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_,
         SUM_0_;
  wire   n1;
  wire   [7:2] carry;

  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(SUM_8_), .S(SUM_7_) );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_add_0 ( A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, 
        B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_9_, SUM_8_, 
        SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_8_, B_7_, B_6_,
         B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_,
         SUM_1_, SUM_0_;
  wire   carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n1;

  ADDFX2 U1_3 ( .A(A_3_), .B(B_3_), .CI(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  ADDFX2 U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFX2 U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  CMPR32X2 U1_8 ( .A(A_8_), .B(B_8_), .C(carry_8_), .CO(SUM_9_), .S(SUM_8_) );
  ADDFX1 U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  ADDFX1 U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module MC2_DW01_inc_2 ( SUM, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_ );
  output [8:0] SUM;
  input A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_;

  wire   [7:2] carry;

  ADDHXL U1_1_2 ( .A(A_2_), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A_1_), .B(A_0_), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A_6_), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A_3_), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_5 ( .A(A_5_), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A_4_), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_7 ( .A(A_7_), .B(carry[7]), .CO(SUM[8]), .S(SUM[7]) );
  CLKINVX1 U1 ( .A(A_0_), .Y(SUM[0]) );
endmodule


module MC2 ( CLK, RESET, in, in_valid, out, out_valid );
  input [7:0] in;
  output [8:0] out;
  input CLK, RESET, in_valid;
  output out_valid;
  wire   n3113, finish, N149, N150, N151, N152, N153, N154, N155, N156,
         start_1_, N182, N183, m43_7_, m55_7_, s1, s2, s3, s4, N833, N834,
         N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845,
         N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856,
         N858, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880,
         N881, N882, N883, N885, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N912, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N931, N932, N933, N934, N935, N937, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N999, N1001, N1002, N1003, N1004, N1005,
         N1006, N1007, N1008, a3_8_, a4_8_, a5_8_, a6_8_, N1073, N1074, N1075,
         N1076, N1077, N1078, N1079, N1080, N1291, N1292, N1293, N1294, N1295,
         N1296, N1297, N1298, N1310, N1311, N1312, N1313, N1314, N1315, N1316,
         N1317, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1348,
         N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1402, N1403, N1404,
         N1405, N1406, N1407, N1408, N1409, N1410, n383, n385, n386, n388,
         n390, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n735,
         n736, n737, n738, n739, n740, n741, n742, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n763, n764, n765, n766, n767, n768, n769, n770, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n8330, n1443, n1445, n1448, n1450, n1452, n1454,
         n1456, n1458, n1459, n1461, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1471, n1475, n1476, n1477, n1478, n1479, n1481, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, N956, N955, N954,
         N953, N952, N951, N950, N949, N948, N986, N985, N984, N983, N982,
         N981, N980, N979, N978, sub_404_carry_2_, sub_404_carry_3_,
         sub_404_carry_4_, sub_404_carry_5_, sub_404_carry_6_,
         sub_404_carry_7_, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1892, n1894, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1969, n1970, n2087, n2088,
         n2089, n2090, n2091, n2092, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108;
  wire   [7:0] mode;
  wire   [7:0] c11;
  wire   [7:0] c12;
  wire   [7:0] c21;
  wire   [7:0] c22;
  wire   [7:0] t11;
  wire   [7:1] t21;
  wire   [7:0] t12;
  wire   [7:0] t22;
  wire   [7:0] node;
  wire   [7:1] max11;
  wire   [7:1] max12;
  wire   [7:1] max21;
  wire   [7:1] max22;
  wire   [8:0] a2;
  wire   [1:0] a1;
  wire   [7:0] outmode;
  wire   [7:2] sub_522_S2_carry;
  wire   [7:2] sub_520_S2_carry;
  wire   [7:2] sub_518_S2_carry;
  wire   [7:2] sub_516_S2_carry;

  MC2_DW01_inc_0 add_439 ( .A(outmode), .SUM({N1080, N1079, N1078, N1077, 
        N1076, N1075, N1074, N1073}) );
  MC2_DW01_sub_5 sub_397 ( .A(t22), .B(c22), .DIFF({N929, N928, N927, N926, 
        N925, N924, N923, N922}) );
  MC2_DW01_sub_6 sub_392 ( .A(c22), .B(t22), .DIFF({N921, N920, N919, N918, 
        N917, N916, N915, N914}) );
  MC2_DW01_sub_7 sub_386 ( .A({t21, n1898}), .B(c21), .DIFF({N902, N901, N900, 
        N899, N898, N897, N896, N895}) );
  MC2_DW01_sub_8 sub_381 ( .A(c21), .B({t21, n1898}), .DIFF({N894, N893, N892, 
        N891, N890, N889, N888, N887}) );
  MC2_DW01_sub_9 sub_375 ( .A(t12), .B(c12), .DIFF({N875, N874, N873, N872, 
        N871, N870, N869, N868}) );
  MC2_DW01_sub_10 sub_370 ( .A(c12), .B(t12), .DIFF({N867, N866, N865, N864, 
        N863, N862, N861, N860}) );
  MC2_DW01_sub_11 sub_364 ( .A(t11), .B(c11), .DIFF({N848, N847, N846, N845, 
        N844, N843, N842, N841}) );
  MC2_DW01_sub_12 sub_359 ( .A(c11), .B(t11), .DIFF({N840, N839, N838, N837, 
        N836, N835, N834, N833}) );
  MC2_DW01_inc_1 r570 ( .A({mode[7], n2785, mode[5:0]}), .SUM({N156, N155, 
        N154, N153, N152, N151, N150, N149}) );
  MC2_DW01_add_5 add_1_root_add_0_root_add_400_3 ( .A_7_(N883), .A_6_(N882), 
        .A_5_(N881), .A_4_(N880), .A_3_(N879), .A_2_(N878), .A_1_(N877), 
        .A_0_(N876), .B_7_(N937), .B_6_(n1917), .B_5_(N935), .B_4_(N934), 
        .B_3_(N933), .B_2_(N932), .B_1_(N931), .B_0_(n1942), .SUM_8_(n3108), 
        .SUM_7_(n3107), .SUM_6_(n3106), .SUM_5_(n3105), .SUM_4_(n3104), 
        .SUM_3_(n3103), .SUM_2_(n3102), .SUM_1_(n3101), .SUM_0_(n3100) );
  MC2_DW01_add_4 add_2_root_add_0_root_add_400_3 ( .A_7_(N856), .A_6_(N855), 
        .A_5_(N854), .A_4_(N853), .A_3_(N852), .A_2_(N851), .A_1_(N850), 
        .A_0_(N849), .B_7_(N910), .B_6_(N909), .B_5_(N908), .B_4_(N907), 
        .B_3_(N906), .B_2_(N905), .B_1_(N904), .B_0_(N903), .SUM_8_(N956), 
        .SUM_7_(N955), .SUM_6_(N954), .SUM_5_(N953), .SUM_4_(N952), .SUM_3_(
        N951), .SUM_2_(N950), .SUM_1_(N949), .SUM_0_(N948) );
  MC2_DW01_add_3 add_0_root_add_0_root_add_400_3 ( .A_8_(N956), .A_7_(N955), 
        .A_6_(N954), .A_5_(N953), .A_4_(N952), .A_3_(N951), .A_2_(N950), 
        .A_1_(N949), .A_0_(N948), .B_8_(n3108), .B_7_(n3107), .B_6_(n3106), 
        .B_5_(n3105), .B_4_(n3104), .B_3_(n3103), .B_2_(n3102), .B_1_(n3101), 
        .B_0_(n3100), .SUM_9_(N967), .SUM_8_(N966), .SUM_7_(N965), .SUM_6_(
        N964), .SUM_5_(N963), .SUM_4_(N962), .SUM_3_(N961), .SUM_2_(N960), 
        .SUM_1_(N959), .SUM_0_(N958) );
  MC2_DW01_add_2 add_1_root_r590 ( .A_7_(max21[7]), .A_6_(max21[6]), .A_5_(
        max21[5]), .A_4_(max21[4]), .A_3_(max21[3]), .A_2_(max21[2]), .A_1_(
        max21[1]), .A_0_(N1329), .B_7_(max22[7]), .B_6_(max22[6]), .B_5_(
        max22[5]), .B_4_(max22[4]), .B_3_(max22[3]), .B_2_(max22[2]), .B_1_(
        max22[1]), .B_0_(N1348), .SUM_8_(n3094), .SUM_7_(n3093), .SUM_6_(n3092), .SUM_5_(n3091), .SUM_4_(n3090), .SUM_3_(n3089), .SUM_2_(n3088), .SUM_1_(
        n3087), .SUM_0_(n3086) );
  MC2_DW01_add_1 add_2_root_r590 ( .A_7_(max11[7]), .A_6_(max11[6]), .A_5_(
        max11[5]), .A_4_(max11[4]), .A_3_(max11[3]), .A_2_(max11[2]), .A_1_(
        max11[1]), .A_0_(N1291), .B_7_(max12[7]), .B_6_(max12[6]), .B_5_(
        max12[5]), .B_4_(max12[4]), .B_3_(max12[3]), .B_2_(max12[2]), .B_1_(
        max12[1]), .B_0_(N1310), .SUM_8_(N986), .SUM_7_(N985), .SUM_6_(N984), 
        .SUM_5_(N983), .SUM_4_(N982), .SUM_3_(N981), .SUM_2_(N980), .SUM_1_(
        N979), .SUM_0_(N978) );
  MC2_DW01_add_0 add_0_root_r590 ( .A_8_(N986), .A_7_(N985), .A_6_(N984), 
        .A_5_(N983), .A_4_(N982), .A_3_(N981), .A_2_(N980), .A_1_(N979), 
        .A_0_(N978), .B_8_(n3094), .B_7_(n3093), .B_6_(n3092), .B_5_(n3091), 
        .B_4_(n3090), .B_3_(n3089), .B_2_(n3088), .B_1_(n3087), .B_0_(n3086), 
        .SUM_9_(N997), .SUM_8_(N996), .SUM_7_(N995), .SUM_6_(N994), .SUM_5_(
        N993), .SUM_4_(N992), .SUM_3_(N991), .SUM_2_(N990), .SUM_1_(N989), 
        .SUM_0_(N988) );
  MC2_DW01_inc_2 add_524_S2_4 ( .SUM({N1410, N1409, N1408, N1407, N1406, N1405, 
        N1404, N1403, N1402}), .A_7_(N997), .A_6_(N996), .A_5_(N995), .A_4_(
        N994), .A_3_(N993), .A_2_(N992), .A_1_(N991), .A_0_(N990) );
  EDFFXL m51_reg_0_ ( .D(n2168), .E(n1464), .CK(CLK), .QN(n640) );
  DFFQX1 a2_reg_8_ ( .D(n1562), .CK(CLK), .Q(a2[8]) );
  DFFQX1 a2_reg_7_ ( .D(n1563), .CK(CLK), .Q(a2[7]) );
  DFFQX1 a2_reg_6_ ( .D(n1564), .CK(CLK), .Q(a2[6]) );
  DFFQX1 a2_reg_5_ ( .D(n1565), .CK(CLK), .Q(a2[5]) );
  DFFQX1 a2_reg_4_ ( .D(n1566), .CK(CLK), .Q(a2[4]) );
  DFFQX1 a2_reg_3_ ( .D(n1567), .CK(CLK), .Q(a2[3]) );
  DFFQX1 a2_reg_2_ ( .D(n1568), .CK(CLK), .Q(a2[2]) );
  EDFFX1 m11_reg_7_ ( .D(n2155), .E(n1838), .CK(CLK), .QN(n441) );
  EDFFX1 m11_reg_6_ ( .D(n2156), .E(n1838), .CK(CLK), .QN(n442) );
  EDFFX1 m11_reg_5_ ( .D(n2158), .E(n1838), .CK(CLK), .QN(n443) );
  EDFFX1 m11_reg_4_ ( .D(n2160), .E(n1838), .CK(CLK), .QN(n444) );
  EDFFX1 m11_reg_3_ ( .D(n2162), .E(n1838), .CK(CLK), .QN(n445) );
  EDFFX1 m11_reg_2_ ( .D(n2164), .E(n1838), .CK(CLK), .QN(n446) );
  EDFFX1 m11_reg_1_ ( .D(n2166), .E(n1838), .CK(CLK), .QN(n447) );
  EDFFX1 m11_reg_0_ ( .D(n2169), .E(n1838), .CK(CLK), .QN(n448) );
  DFFQX1 a6_reg_8_ ( .D(n1526), .CK(CLK), .Q(a6_8_) );
  EDFFX1 m16_reg_7_ ( .D(n2155), .E(n1487), .CK(CLK), .QN(n481) );
  EDFFX1 m16_reg_6_ ( .D(n2157), .E(n1487), .CK(CLK), .QN(n482) );
  EDFFX1 m16_reg_5_ ( .D(n2159), .E(n1487), .CK(CLK), .QN(n483) );
  EDFFX1 m16_reg_4_ ( .D(n2161), .E(n1487), .CK(CLK), .QN(n484) );
  EDFFX1 m16_reg_3_ ( .D(n2163), .E(n1487), .CK(CLK), .QN(n485) );
  EDFFX1 m16_reg_2_ ( .D(n2165), .E(n1487), .CK(CLK), .QN(n486) );
  EDFFX1 m16_reg_1_ ( .D(n2167), .E(n1487), .CK(CLK), .QN(n487) );
  EDFFX1 m16_reg_0_ ( .D(n2168), .E(n1487), .CK(CLK), .QN(n488) );
  EDFFX1 m61_reg_7_ ( .D(n2154), .E(n1454), .CK(CLK), .QN(n2314) );
  EDFFX1 m66_reg_7_ ( .D(n2154), .E(n1443), .CK(CLK), .QN(n2313) );
  DFFQX1 a5_reg_8_ ( .D(n1535), .CK(CLK), .Q(a5_8_) );
  DFFQX1 a4_reg_8_ ( .D(n1544), .CK(CLK), .Q(a4_8_) );
  DFFQX1 a3_reg_8_ ( .D(n1553), .CK(CLK), .Q(a3_8_) );
  EDFFX1 m14_reg_7_ ( .D(n2154), .E(n1489), .CK(CLK), .QN(n465) );
  EDFFX1 m14_reg_6_ ( .D(n2156), .E(n1489), .CK(CLK), .QN(n466) );
  EDFFX1 m14_reg_5_ ( .D(n2158), .E(n1489), .CK(CLK), .QN(n467) );
  EDFFX1 m14_reg_4_ ( .D(n2160), .E(n1489), .CK(CLK), .QN(n468) );
  EDFFX1 m14_reg_3_ ( .D(n2162), .E(n1489), .CK(CLK), .QN(n469) );
  EDFFX1 m14_reg_2_ ( .D(n2164), .E(n1489), .CK(CLK), .QN(n470) );
  EDFFX1 m14_reg_1_ ( .D(n2166), .E(n1489), .CK(CLK), .QN(n471) );
  EDFFX1 m14_reg_0_ ( .D(n2168), .E(n1489), .CK(CLK), .QN(n472) );
  EDFFX1 m13_reg_7_ ( .D(n2155), .E(n1490), .CK(CLK), .QN(n457) );
  EDFFX1 m12_reg_7_ ( .D(n2155), .E(n1839), .CK(CLK), .QN(n449) );
  EDFFX1 m12_reg_6_ ( .D(n2157), .E(n1839), .CK(CLK), .QN(n450) );
  EDFFX1 m12_reg_5_ ( .D(n2159), .E(n1839), .CK(CLK), .QN(n451) );
  EDFFX1 m12_reg_4_ ( .D(n2161), .E(n1839), .CK(CLK), .QN(n452) );
  EDFFX1 m12_reg_3_ ( .D(n2163), .E(n1839), .CK(CLK), .QN(n453) );
  EDFFX1 m12_reg_2_ ( .D(n2165), .E(n1839), .CK(CLK), .QN(n454) );
  EDFFX1 m12_reg_1_ ( .D(n2167), .E(n1839), .CK(CLK), .QN(n455) );
  EDFFX1 m12_reg_0_ ( .D(n2169), .E(n1839), .CK(CLK), .QN(n456) );
  EDFFX1 m15_reg_7_ ( .D(n3076), .E(n1488), .CK(CLK), .QN(n473) );
  EDFFX1 m15_reg_6_ ( .D(n2157), .E(n1488), .CK(CLK), .QN(n474) );
  EDFFX1 m15_reg_5_ ( .D(n2159), .E(n1488), .CK(CLK), .QN(n475) );
  EDFFX1 m15_reg_4_ ( .D(n2161), .E(n1488), .CK(CLK), .QN(n476) );
  EDFFX1 m15_reg_3_ ( .D(n2163), .E(n1488), .CK(CLK), .QN(n477) );
  EDFFX1 m15_reg_2_ ( .D(n2165), .E(n1488), .CK(CLK), .QN(n478) );
  EDFFX1 m15_reg_1_ ( .D(n2167), .E(n1488), .CK(CLK), .QN(n479) );
  EDFFX1 m15_reg_0_ ( .D(n2169), .E(n1488), .CK(CLK), .QN(n480) );
  EDFFX1 m21_reg_7_ ( .D(n2154), .E(n1486), .CK(CLK), .QN(n489) );
  EDFFX1 m21_reg_6_ ( .D(n2156), .E(n1486), .CK(CLK), .QN(n490) );
  EDFFX1 m21_reg_5_ ( .D(n2158), .E(n1486), .CK(CLK), .QN(n491) );
  EDFFX1 m21_reg_4_ ( .D(n2160), .E(n1486), .CK(CLK), .QN(n492) );
  EDFFX1 m21_reg_3_ ( .D(n2162), .E(n1486), .CK(CLK), .QN(n493) );
  EDFFX1 m21_reg_2_ ( .D(n2164), .E(n1486), .CK(CLK), .QN(n494) );
  EDFFX1 m21_reg_1_ ( .D(n2166), .E(n1486), .CK(CLK), .QN(n495) );
  EDFFX1 m21_reg_0_ ( .D(n2168), .E(n1486), .CK(CLK), .QN(n496) );
  EDFFX1 m62_reg_7_ ( .D(n2154), .E(n1452), .CK(CLK), .QN(n422) );
  EDFFX1 m46_reg_7_ ( .D(n2155), .E(n1465), .CK(CLK), .QN(n625) );
  EDFFX1 m46_reg_6_ ( .D(n2157), .E(n1465), .CK(CLK), .QN(n626) );
  EDFFX1 m46_reg_5_ ( .D(n2159), .E(n1465), .CK(CLK), .QN(n627) );
  EDFFX1 m46_reg_4_ ( .D(n2161), .E(n1465), .CK(CLK), .QN(n628) );
  EDFFX1 m46_reg_3_ ( .D(n2163), .E(n1465), .CK(CLK), .QN(n629) );
  EDFFX1 m46_reg_2_ ( .D(n2165), .E(n1465), .CK(CLK), .QN(n630) );
  EDFFX1 m46_reg_1_ ( .D(n2167), .E(n1465), .CK(CLK), .QN(n631) );
  EDFFX1 m46_reg_0_ ( .D(n2169), .E(n1465), .CK(CLK), .QN(n632) );
  EDFFX1 m56_reg_7_ ( .D(n2155), .E(n1456), .CK(CLK), .QN(n673) );
  EDFFX1 m65_reg_7_ ( .D(n2155), .E(n1445), .CK(CLK), .QN(n2315) );
  EDFFX1 m51_reg_7_ ( .D(n2155), .E(n1464), .CK(CLK), .QN(n633) );
  EDFFX1 m51_reg_6_ ( .D(n3077), .E(n1464), .CK(CLK), .QN(n634) );
  EDFFX1 m51_reg_5_ ( .D(n2159), .E(n1464), .CK(CLK), .QN(n635) );
  EDFFX1 m51_reg_4_ ( .D(n2161), .E(n1464), .CK(CLK), .QN(n636) );
  EDFFX1 m51_reg_3_ ( .D(n3080), .E(n1464), .CK(CLK), .QN(n637) );
  EDFFX1 m51_reg_2_ ( .D(n2165), .E(n1464), .CK(CLK), .QN(n638) );
  EDFFX1 m51_reg_1_ ( .D(n3082), .E(n1464), .CK(CLK), .QN(n639) );
  EDFFX1 m36_reg_7_ ( .D(n2155), .E(n1841), .CK(CLK), .Q(n1821), .QN(n577) );
  EDFFX1 m36_reg_6_ ( .D(n2157), .E(n1841), .CK(CLK), .Q(n1820), .QN(n578) );
  EDFFX1 m36_reg_5_ ( .D(n2159), .E(n1841), .CK(CLK), .Q(n1819), .QN(n579) );
  EDFFX1 m36_reg_4_ ( .D(n2161), .E(n1841), .CK(CLK), .Q(n1818), .QN(n580) );
  EDFFX1 m36_reg_3_ ( .D(n2163), .E(n1841), .CK(CLK), .Q(n1817), .QN(n581) );
  EDFFX1 m36_reg_2_ ( .D(n2165), .E(n1841), .CK(CLK), .Q(n1816), .QN(n582) );
  EDFFX1 m36_reg_1_ ( .D(n2167), .E(n1841), .CK(CLK), .Q(n1815), .QN(n583) );
  EDFFX1 m36_reg_0_ ( .D(n2169), .E(n1841), .CK(CLK), .Q(n1814), .QN(n584) );
  EDFFX1 m26_reg_7_ ( .D(n2154), .E(n1479), .CK(CLK), .Q(n1813), .QN(n529) );
  EDFFX1 m26_reg_6_ ( .D(n2156), .E(n1479), .CK(CLK), .Q(n1812), .QN(n530) );
  EDFFX1 m26_reg_5_ ( .D(n2158), .E(n1479), .CK(CLK), .Q(n1811), .QN(n531) );
  EDFFX1 m26_reg_4_ ( .D(n2160), .E(n1479), .CK(CLK), .Q(n1810), .QN(n532) );
  EDFFX1 m26_reg_3_ ( .D(n2162), .E(n1479), .CK(CLK), .Q(n1809), .QN(n533) );
  EDFFX1 m26_reg_2_ ( .D(n2164), .E(n1479), .CK(CLK), .Q(n1808), .QN(n534) );
  EDFFX1 m26_reg_1_ ( .D(n2166), .E(n1479), .CK(CLK), .Q(n1807), .QN(n535) );
  EDFFX1 m26_reg_0_ ( .D(n2168), .E(n1479), .CK(CLK), .Q(n1806), .QN(n536) );
  EDFFX1 m63_reg_7_ ( .D(n2155), .E(n1450), .CK(CLK), .Q(n1773), .QN(n399) );
  EDFFX1 m64_reg_7_ ( .D(n2155), .E(n1448), .CK(CLK), .Q(n1805), .QN(n407) );
  EDFFX1 m64_reg_6_ ( .D(n2157), .E(n1448), .CK(CLK), .Q(n1804), .QN(n408) );
  EDFFX1 m64_reg_5_ ( .D(n2159), .E(n1448), .CK(CLK), .Q(n1803), .QN(n409) );
  EDFFX1 m64_reg_4_ ( .D(n2161), .E(n1448), .CK(CLK), .Q(n1802), .QN(n410) );
  EDFFX1 m64_reg_3_ ( .D(n2163), .E(n1448), .CK(CLK), .Q(n1801), .QN(n411) );
  EDFFX1 m64_reg_2_ ( .D(n2165), .E(n1448), .CK(CLK), .Q(n1800), .QN(n412) );
  EDFFX1 m64_reg_1_ ( .D(n2167), .E(n1448), .CK(CLK), .Q(n1799), .QN(n413) );
  EDFFX1 m64_reg_0_ ( .D(n2169), .E(n1448), .CK(CLK), .Q(n1798), .QN(n414) );
  DFFQX1 a1_reg_0_ ( .D(n1516), .CK(CLK), .Q(a1[0]) );
  DFFQX1 a2_reg_0_ ( .D(n3072), .CK(CLK), .Q(a2[0]) );
  DFFQX1 a2_reg_1_ ( .D(n1569), .CK(CLK), .Q(a2[1]) );
  EDFFX1 m22_reg_7_ ( .D(n2155), .E(n1485), .CK(CLK), .QN(n497) );
  EDFFX1 m22_reg_6_ ( .D(n2157), .E(n1485), .CK(CLK), .QN(n498) );
  EDFFX1 m22_reg_5_ ( .D(n2159), .E(n1485), .CK(CLK), .QN(n499) );
  EDFFX1 m22_reg_4_ ( .D(n2161), .E(n1485), .CK(CLK), .QN(n500) );
  EDFFX1 m22_reg_3_ ( .D(n2163), .E(n1485), .CK(CLK), .QN(n501) );
  EDFFX1 m22_reg_2_ ( .D(n2165), .E(n1485), .CK(CLK), .QN(n502) );
  EDFFX1 m22_reg_1_ ( .D(n2167), .E(n1485), .CK(CLK), .QN(n503) );
  EDFFX1 m22_reg_0_ ( .D(n2169), .E(n1485), .CK(CLK), .QN(n504) );
  EDFFX1 m52_reg_7_ ( .D(n2155), .E(n1463), .CK(CLK), .QN(n641) );
  EDFFX1 m52_reg_6_ ( .D(n2157), .E(n1463), .CK(CLK), .QN(n642) );
  EDFFX1 m52_reg_5_ ( .D(n2159), .E(n1463), .CK(CLK), .QN(n643) );
  EDFFX1 m52_reg_4_ ( .D(n2161), .E(n1463), .CK(CLK), .QN(n644) );
  EDFFX1 m52_reg_3_ ( .D(n2163), .E(n1463), .CK(CLK), .QN(n645) );
  EDFFX1 m52_reg_2_ ( .D(n2165), .E(n1463), .CK(CLK), .QN(n646) );
  EDFFX1 m52_reg_1_ ( .D(n2167), .E(n1463), .CK(CLK), .QN(n647) );
  EDFFX1 m52_reg_0_ ( .D(n2169), .E(n1463), .CK(CLK), .QN(n648) );
  EDFFX1 m44_reg_7_ ( .D(n2155), .E(n1467), .CK(CLK), .QN(n609) );
  EDFFX1 m44_reg_6_ ( .D(n3077), .E(n1467), .CK(CLK), .QN(n610) );
  EDFFX1 m44_reg_5_ ( .D(n3078), .E(n1467), .CK(CLK), .QN(n611) );
  EDFFX1 m44_reg_4_ ( .D(n3079), .E(n1467), .CK(CLK), .QN(n612) );
  EDFFX1 m44_reg_3_ ( .D(n3080), .E(n1467), .CK(CLK), .QN(n613) );
  EDFFX1 m44_reg_2_ ( .D(n3081), .E(n1467), .CK(CLK), .QN(n614) );
  EDFFX1 m44_reg_1_ ( .D(n3082), .E(n1467), .CK(CLK), .QN(n615) );
  EDFFX1 m44_reg_0_ ( .D(n3083), .E(n1467), .CK(CLK), .QN(n616) );
  EDFFX1 m45_reg_7_ ( .D(n2154), .E(n1466), .CK(CLK), .QN(n617) );
  EDFFX1 m45_reg_6_ ( .D(n2156), .E(n1466), .CK(CLK), .QN(n618) );
  EDFFX1 m45_reg_5_ ( .D(n2158), .E(n1466), .CK(CLK), .QN(n619) );
  EDFFX1 m45_reg_4_ ( .D(n2160), .E(n1466), .CK(CLK), .QN(n620) );
  EDFFX1 m45_reg_3_ ( .D(n2162), .E(n1466), .CK(CLK), .QN(n621) );
  EDFFX1 m45_reg_2_ ( .D(n2164), .E(n1466), .CK(CLK), .QN(n622) );
  EDFFX1 m45_reg_1_ ( .D(n2166), .E(n1466), .CK(CLK), .QN(n623) );
  EDFFX1 m45_reg_0_ ( .D(n2168), .E(n1466), .CK(CLK), .QN(n624) );
  EDFFX1 m55_reg_6_ ( .D(n2157), .E(n1458), .CK(CLK), .QN(n666) );
  EDFFX1 m55_reg_5_ ( .D(n2159), .E(n1458), .CK(CLK), .QN(n667) );
  EDFFX1 m55_reg_4_ ( .D(n2161), .E(n1458), .CK(CLK), .QN(n668) );
  EDFFX1 m55_reg_3_ ( .D(n2163), .E(n1458), .CK(CLK), .QN(n669) );
  EDFFX1 m55_reg_2_ ( .D(n2165), .E(n1458), .CK(CLK), .QN(n670) );
  EDFFX1 m55_reg_1_ ( .D(n2167), .E(n1458), .CK(CLK), .QN(n671) );
  EDFFX1 m55_reg_0_ ( .D(n2169), .E(n1458), .CK(CLK), .QN(n672) );
  EDFFX1 m53_reg_7_ ( .D(n2155), .E(n1461), .CK(CLK), .Q(n1765), .QN(n649) );
  EDFFX1 m53_reg_6_ ( .D(n3077), .E(n1461), .CK(CLK), .Q(n1764), .QN(n650) );
  EDFFX1 m53_reg_5_ ( .D(n3078), .E(n1461), .CK(CLK), .Q(n1763), .QN(n651) );
  EDFFX1 m53_reg_4_ ( .D(n3079), .E(n1461), .CK(CLK), .Q(n1762), .QN(n652) );
  EDFFX1 m53_reg_3_ ( .D(n3080), .E(n1461), .CK(CLK), .Q(n1761), .QN(n653) );
  EDFFX1 m53_reg_2_ ( .D(n3081), .E(n1461), .CK(CLK), .Q(n1760), .QN(n654) );
  EDFFX1 m53_reg_1_ ( .D(n3082), .E(n1461), .CK(CLK), .Q(n1759), .QN(n655) );
  EDFFX1 m53_reg_0_ ( .D(n3083), .E(n1461), .CK(CLK), .Q(n1758), .QN(n656) );
  EDFFX1 m54_reg_7_ ( .D(n2154), .E(n1459), .CK(CLK), .Q(n1789), .QN(n657) );
  EDFFX1 m54_reg_6_ ( .D(n2156), .E(n1459), .CK(CLK), .Q(n1788), .QN(n658) );
  EDFFX1 m54_reg_5_ ( .D(n2158), .E(n1459), .CK(CLK), .Q(n1787), .QN(n659) );
  EDFFX1 m54_reg_4_ ( .D(n2160), .E(n1459), .CK(CLK), .Q(n1786), .QN(n660) );
  EDFFX1 m54_reg_3_ ( .D(n2162), .E(n1459), .CK(CLK), .Q(n1785), .QN(n661) );
  EDFFX1 m54_reg_2_ ( .D(n2164), .E(n1459), .CK(CLK), .Q(n1784), .QN(n662) );
  EDFFX1 m54_reg_1_ ( .D(n2166), .E(n1459), .CK(CLK), .Q(n1783), .QN(n663) );
  EDFFX1 m54_reg_0_ ( .D(n2168), .E(n1459), .CK(CLK), .Q(n1782), .QN(n664) );
  DFFQX1 m55_reg_7_ ( .D(n1654), .CK(CLK), .Q(m55_7_) );
  DFFQX1 m43_reg_7_ ( .D(n1655), .CK(CLK), .Q(m43_7_) );
  EDFFX1 m31_reg_7_ ( .D(n2155), .E(n1478), .CK(CLK), .Q(n1837), .QN(n537) );
  EDFFX1 m31_reg_6_ ( .D(n2157), .E(n1478), .CK(CLK), .Q(n1836), .QN(n538) );
  EDFFX1 m31_reg_5_ ( .D(n2159), .E(n1478), .CK(CLK), .Q(n1835), .QN(n539) );
  EDFFX1 m31_reg_4_ ( .D(n2161), .E(n1478), .CK(CLK), .Q(n1834), .QN(n540) );
  EDFFX1 m31_reg_3_ ( .D(n2163), .E(n1478), .CK(CLK), .Q(n1833), .QN(n541) );
  EDFFX1 m31_reg_2_ ( .D(n2165), .E(n1478), .CK(CLK), .Q(n1832), .QN(n542) );
  EDFFX1 m31_reg_1_ ( .D(n2167), .E(n1478), .CK(CLK), .Q(n1831), .QN(n543) );
  EDFFX1 m31_reg_0_ ( .D(n2169), .E(n1478), .CK(CLK), .Q(n1830), .QN(n544) );
  EDFFX1 m41_reg_7_ ( .D(n2155), .E(n1471), .CK(CLK), .Q(n1829), .QN(n585) );
  EDFFX1 m41_reg_6_ ( .D(n2156), .E(n1471), .CK(CLK), .Q(n1828), .QN(n586) );
  EDFFX1 m41_reg_5_ ( .D(n2158), .E(n1471), .CK(CLK), .Q(n1827), .QN(n587) );
  EDFFX1 m41_reg_4_ ( .D(n2160), .E(n1471), .CK(CLK), .Q(n1826), .QN(n588) );
  EDFFX1 m41_reg_3_ ( .D(n2162), .E(n1471), .CK(CLK), .Q(n1825), .QN(n589) );
  EDFFX1 m41_reg_2_ ( .D(n2164), .E(n1471), .CK(CLK), .Q(n1824), .QN(n590) );
  EDFFX1 m41_reg_1_ ( .D(n2166), .E(n1471), .CK(CLK), .Q(n1823), .QN(n591) );
  EDFFX1 m41_reg_0_ ( .D(n2169), .E(n1471), .CK(CLK), .Q(n1822), .QN(n592) );
  EDFFX1 m24_reg_7_ ( .D(n2155), .E(n1483), .CK(CLK), .Q(n1757), .QN(n513) );
  EDFFX1 m24_reg_6_ ( .D(n2157), .E(n1483), .CK(CLK), .Q(n1756), .QN(n514) );
  EDFFX1 m24_reg_5_ ( .D(n2159), .E(n1483), .CK(CLK), .Q(n1755), .QN(n515) );
  EDFFX1 m24_reg_4_ ( .D(n2161), .E(n1483), .CK(CLK), .Q(n1754), .QN(n516) );
  EDFFX1 m24_reg_3_ ( .D(n2163), .E(n1483), .CK(CLK), .Q(n1753), .QN(n517) );
  EDFFX1 m24_reg_2_ ( .D(n2165), .E(n1483), .CK(CLK), .Q(n1752), .QN(n518) );
  EDFFX1 m24_reg_1_ ( .D(n2167), .E(n1483), .CK(CLK), .Q(n1751), .QN(n519) );
  EDFFX1 m24_reg_0_ ( .D(n2169), .E(n1483), .CK(CLK), .Q(n1750), .QN(n520) );
  EDFFX1 m25_reg_7_ ( .D(n2155), .E(n1481), .CK(CLK), .Q(n1717), .QN(n521) );
  EDFFX1 m25_reg_6_ ( .D(n2157), .E(n1481), .CK(CLK), .Q(n1716), .QN(n522) );
  EDFFX1 m25_reg_5_ ( .D(n3078), .E(n1481), .CK(CLK), .Q(n1715), .QN(n523) );
  EDFFX1 m25_reg_4_ ( .D(n3079), .E(n1481), .CK(CLK), .Q(n1714), .QN(n524) );
  EDFFX1 m25_reg_3_ ( .D(n2163), .E(n1481), .CK(CLK), .Q(n1713), .QN(n525) );
  EDFFX1 m25_reg_2_ ( .D(n3081), .E(n1481), .CK(CLK), .Q(n1712), .QN(n526) );
  EDFFX1 m25_reg_1_ ( .D(n2167), .E(n1481), .CK(CLK), .Q(n1711), .QN(n527) );
  EDFFX1 m25_reg_0_ ( .D(n3083), .E(n1481), .CK(CLK), .Q(n1710), .QN(n528) );
  EDFFX1 m35_reg_7_ ( .D(n2155), .E(n1840), .CK(CLK), .Q(n1709), .QN(n569) );
  EDFFX1 m35_reg_6_ ( .D(n3077), .E(n1840), .CK(CLK), .Q(n1708), .QN(n570) );
  EDFFX1 m35_reg_5_ ( .D(n3078), .E(n1840), .CK(CLK), .Q(n1707), .QN(n571) );
  EDFFX1 m35_reg_4_ ( .D(n3079), .E(n1840), .CK(CLK), .Q(n1706), .QN(n572) );
  EDFFX1 m35_reg_3_ ( .D(n3080), .E(n1840), .CK(CLK), .Q(n1705), .QN(n573) );
  EDFFX1 m35_reg_2_ ( .D(n3081), .E(n1840), .CK(CLK), .Q(n1704), .QN(n574) );
  EDFFX1 m35_reg_1_ ( .D(n3082), .E(n1840), .CK(CLK), .Q(n1703), .QN(n575) );
  EDFFX1 m35_reg_0_ ( .D(n3083), .E(n1840), .CK(CLK), .Q(n1702), .QN(n576) );
  EDFFX1 m34_reg_7_ ( .D(n2155), .E(n1475), .CK(CLK), .Q(n1749), .QN(n561) );
  EDFFX1 m34_reg_6_ ( .D(n2157), .E(n1475), .CK(CLK), .Q(n1748), .QN(n562) );
  EDFFX1 m34_reg_5_ ( .D(n2159), .E(n1475), .CK(CLK), .Q(n1747), .QN(n563) );
  EDFFX1 m34_reg_4_ ( .D(n2161), .E(n1475), .CK(CLK), .Q(n1746), .QN(n564) );
  EDFFX1 m34_reg_3_ ( .D(n2163), .E(n1475), .CK(CLK), .Q(n1745), .QN(n565) );
  EDFFX1 m34_reg_2_ ( .D(n2165), .E(n1475), .CK(CLK), .Q(n1744), .QN(n566) );
  EDFFX1 m34_reg_1_ ( .D(n2167), .E(n1475), .CK(CLK), .Q(n1743), .QN(n567) );
  EDFFX1 m34_reg_0_ ( .D(n2169), .E(n1475), .CK(CLK), .Q(n1742), .QN(n568) );
  EDFFX1 m32_reg_7_ ( .D(n2155), .E(n1477), .CK(CLK), .Q(n1733), .QN(n545) );
  EDFFX1 m32_reg_6_ ( .D(n3077), .E(n1477), .CK(CLK), .Q(n1732), .QN(n546) );
  EDFFX1 m32_reg_5_ ( .D(n3078), .E(n1477), .CK(CLK), .Q(n1731), .QN(n547) );
  EDFFX1 m32_reg_4_ ( .D(n3079), .E(n1477), .CK(CLK), .Q(n1730), .QN(n548) );
  EDFFX1 m32_reg_3_ ( .D(n3080), .E(n1477), .CK(CLK), .Q(n1729), .QN(n549) );
  EDFFX1 m32_reg_2_ ( .D(n3081), .E(n1477), .CK(CLK), .Q(n1728), .QN(n550) );
  EDFFX1 m32_reg_1_ ( .D(n3082), .E(n1477), .CK(CLK), .Q(n1727), .QN(n551) );
  EDFFX1 m32_reg_0_ ( .D(n3083), .E(n1477), .CK(CLK), .Q(n1726), .QN(n552) );
  EDFFX1 m42_reg_7_ ( .D(n2154), .E(n1469), .CK(CLK), .Q(n1725), .QN(n593) );
  EDFFX1 m42_reg_6_ ( .D(n2156), .E(n1469), .CK(CLK), .Q(n1724), .QN(n594) );
  EDFFX1 m42_reg_5_ ( .D(n2158), .E(n1469), .CK(CLK), .Q(n1723), .QN(n595) );
  EDFFX1 m42_reg_4_ ( .D(n2160), .E(n1469), .CK(CLK), .Q(n1722), .QN(n596) );
  EDFFX1 m42_reg_3_ ( .D(n2162), .E(n1469), .CK(CLK), .Q(n1721), .QN(n597) );
  EDFFX1 m42_reg_2_ ( .D(n2164), .E(n1469), .CK(CLK), .Q(n1720), .QN(n598) );
  EDFFX1 m42_reg_1_ ( .D(n2166), .E(n1469), .CK(CLK), .Q(n1719), .QN(n599) );
  EDFFX1 m42_reg_0_ ( .D(n2168), .E(n1469), .CK(CLK), .Q(n1718), .QN(n600) );
  EDFFX1 m33_reg_7_ ( .D(n2154), .E(n1476), .CK(CLK), .Q(n1696), .QN(n553) );
  EDFFX1 m33_reg_6_ ( .D(n2156), .E(n1476), .CK(CLK), .Q(n1695), .QN(n554) );
  EDFFX1 m33_reg_5_ ( .D(n2158), .E(n1476), .CK(CLK), .Q(n1694), .QN(n555) );
  EDFFX1 m33_reg_4_ ( .D(n2160), .E(n1476), .CK(CLK), .Q(n1693), .QN(n556) );
  EDFFX1 m33_reg_3_ ( .D(n2162), .E(n1476), .CK(CLK), .Q(n1692), .QN(n557) );
  EDFFX1 m33_reg_2_ ( .D(n2164), .E(n1476), .CK(CLK), .Q(n1691), .QN(n558) );
  EDFFX1 m33_reg_1_ ( .D(n2166), .E(n1476), .CK(CLK), .Q(n1690), .QN(n559) );
  EDFFX1 m33_reg_0_ ( .D(n2168), .E(n1476), .CK(CLK), .Q(n1689), .QN(n560) );
  DFFQX1 a1_reg_1_ ( .D(n1515), .CK(CLK), .Q(a1[1]) );
  EDFFX1 m23_reg_7_ ( .D(n2155), .E(n1484), .CK(CLK), .Q(n1797), .QN(n505) );
  EDFFX1 m23_reg_6_ ( .D(n2157), .E(n1484), .CK(CLK), .Q(n1796), .QN(n506) );
  EDFFX1 m23_reg_5_ ( .D(n2159), .E(n1484), .CK(CLK), .Q(n1795), .QN(n507) );
  EDFFX1 m23_reg_4_ ( .D(n2161), .E(n1484), .CK(CLK), .Q(n1794), .QN(n508) );
  EDFFX1 m23_reg_3_ ( .D(n2163), .E(n1484), .CK(CLK), .Q(n1793), .QN(n509) );
  EDFFX1 m23_reg_2_ ( .D(n2165), .E(n1484), .CK(CLK), .Q(n1792), .QN(n510) );
  EDFFX1 m23_reg_1_ ( .D(n2167), .E(n1484), .CK(CLK), .Q(n1791), .QN(n511) );
  EDFFX1 m23_reg_0_ ( .D(n2169), .E(n1484), .CK(CLK), .Q(n1790), .QN(n512) );
  EDFFX1 m43_reg_6_ ( .D(n2157), .E(n1468), .CK(CLK), .Q(n1772), .QN(n602) );
  EDFFX1 m43_reg_5_ ( .D(n2159), .E(n1468), .CK(CLK), .Q(n1771), .QN(n603) );
  EDFFX1 m43_reg_4_ ( .D(n2161), .E(n1468), .CK(CLK), .Q(n1770), .QN(n604) );
  EDFFX1 m43_reg_3_ ( .D(n2163), .E(n1468), .CK(CLK), .Q(n1769), .QN(n605) );
  EDFFX1 m43_reg_2_ ( .D(n2165), .E(n1468), .CK(CLK), .Q(n1768), .QN(n606) );
  EDFFX1 m43_reg_1_ ( .D(n2167), .E(n1468), .CK(CLK), .Q(n1767), .QN(n607) );
  EDFFX1 m43_reg_0_ ( .D(n2169), .E(n1468), .CK(CLK), .Q(n1766), .QN(n608) );
  EDFFTRX1 outmode_reg_7_ ( .RN(n2170), .D(N1080), .E(n2094), .CK(CLK), .Q(
        outmode[7]) );
  EDFFTRX1 outmode_reg_6_ ( .RN(n2170), .D(N1079), .E(n2094), .CK(CLK), .Q(
        outmode[6]) );
  EDFFTRX1 outmode_reg_5_ ( .RN(n2170), .D(N1078), .E(n2094), .CK(CLK), .Q(
        outmode[5]) );
  EDFFTRX1 outmode_reg_4_ ( .RN(n2170), .D(N1077), .E(n2094), .CK(CLK), .Q(
        outmode[4]) );
  EDFFTRX1 outmode_reg_3_ ( .RN(n2170), .D(N1076), .E(n2094), .CK(CLK), .Q(
        outmode[3]) );
  EDFFTRX1 outmode_reg_2_ ( .RN(n2170), .D(N1075), .E(n2094), .CK(CLK), .Q(
        outmode[2]) );
  EDFFTRX1 outmode_reg_1_ ( .RN(n2170), .D(N1074), .E(n2094), .CK(CLK), .Q(
        outmode[1]) );
  DFFQX1 max21_reg_7_ ( .D(n1582), .CK(CLK), .Q(max21[7]) );
  DFFQX1 max21_reg_6_ ( .D(n1583), .CK(CLK), .Q(max21[6]) );
  DFFQX1 max11_reg_7_ ( .D(n1598), .CK(CLK), .Q(max11[7]) );
  DFFQX1 max11_reg_6_ ( .D(n1599), .CK(CLK), .Q(max11[6]) );
  DFFQX1 max22_reg_6_ ( .D(n1575), .CK(CLK), .Q(max22[6]) );
  DFFQX1 max12_reg_7_ ( .D(n1590), .CK(CLK), .Q(max12[7]) );
  DFFQX1 max12_reg_6_ ( .D(n1591), .CK(CLK), .Q(max12[6]) );
  DFFQX2 node_reg_0_ ( .D(n1613), .CK(CLK), .Q(node[0]) );
  DFFQX1 finish_reg ( .D(n1680), .CK(CLK), .Q(finish) );
  DFFQX2 node_reg_2_ ( .D(n1611), .CK(CLK), .Q(node[2]) );
  DFFQX1 out_valid_reg ( .D(n1681), .CK(CLK), .Q(n3113) );
  DFFQX1 max21_reg_5_ ( .D(n1584), .CK(CLK), .Q(max21[5]) );
  DFFQX1 max21_reg_4_ ( .D(n1585), .CK(CLK), .Q(max21[4]) );
  DFFQX1 max21_reg_3_ ( .D(n1586), .CK(CLK), .Q(max21[3]) );
  DFFQX1 max21_reg_2_ ( .D(n1587), .CK(CLK), .Q(max21[2]) );
  DFFQX1 max11_reg_5_ ( .D(n1600), .CK(CLK), .Q(max11[5]) );
  DFFQX1 max11_reg_4_ ( .D(n1601), .CK(CLK), .Q(max11[4]) );
  DFFQX1 max11_reg_3_ ( .D(n1602), .CK(CLK), .Q(max11[3]) );
  DFFQX1 max11_reg_2_ ( .D(n1603), .CK(CLK), .Q(max11[2]) );
  DFFQX1 node_reg_3_ ( .D(n1610), .CK(CLK), .Q(node[3]) );
  DFFQX1 node_reg_1_ ( .D(n1612), .CK(CLK), .Q(node[1]) );
  DFFQX1 max11_reg_1_ ( .D(n1604), .CK(CLK), .Q(max11[1]) );
  DFFQX1 max21_reg_1_ ( .D(n1588), .CK(CLK), .Q(max21[1]) );
  DFFQX1 max22_reg_5_ ( .D(n1576), .CK(CLK), .Q(max22[5]) );
  DFFQX1 max22_reg_4_ ( .D(n1577), .CK(CLK), .Q(max22[4]) );
  DFFQX1 max22_reg_3_ ( .D(n1578), .CK(CLK), .Q(max22[3]) );
  DFFQX1 max22_reg_2_ ( .D(n1579), .CK(CLK), .Q(max22[2]) );
  DFFQX1 max22_reg_1_ ( .D(n1580), .CK(CLK), .Q(max22[1]) );
  DFFQX1 max12_reg_5_ ( .D(n1592), .CK(CLK), .Q(max12[5]) );
  DFFQX1 max12_reg_4_ ( .D(n1593), .CK(CLK), .Q(max12[4]) );
  DFFQX1 max12_reg_3_ ( .D(n1594), .CK(CLK), .Q(max12[3]) );
  DFFQX1 max12_reg_2_ ( .D(n1595), .CK(CLK), .Q(max12[2]) );
  DFFQX1 c11_reg_7_ ( .D(n1646), .CK(CLK), .Q(c11[7]) );
  DFFQX1 c21_reg_5_ ( .D(n1666), .CK(CLK), .Q(c21[5]) );
  DFFQX1 c11_reg_5_ ( .D(n1648), .CK(CLK), .Q(c11[5]) );
  DFFQX1 c11_reg_3_ ( .D(n1650), .CK(CLK), .Q(c11[3]) );
  DFFQX1 c11_reg_1_ ( .D(n1652), .CK(CLK), .Q(c11[1]) );
  EDFFTRX1 outmode_reg_0_ ( .RN(n2171), .D(N1073), .E(n2094), .CK(CLK), .Q(
        outmode[0]) );
  DFFQX1 max12_reg_1_ ( .D(n1596), .CK(CLK), .Q(max12[1]) );
  DFFQX1 c21_reg_7_ ( .D(n1664), .CK(CLK), .Q(c21[7]) );
  DFFQX1 t21_reg_7_ ( .D(n1638), .CK(CLK), .Q(t21[7]) );
  DFFQX1 c22_reg_5_ ( .D(n1658), .CK(CLK), .Q(c22[5]) );
  DFFQXL s4_reg ( .D(n1570), .CK(CLK), .Q(s4) );
  DFFQXL s3_reg ( .D(n1571), .CK(CLK), .Q(s3) );
  DFFQXL s2_reg ( .D(n1572), .CK(CLK), .Q(s2) );
  DFFQXL node_reg_6_ ( .D(n1607), .CK(CLK), .Q(node[6]) );
  DFFQXL node_reg_5_ ( .D(n1608), .CK(CLK), .Q(node[5]) );
  DFFQXL node_reg_7_ ( .D(n1606), .CK(CLK), .Q(node[7]) );
  DFFQXL node_reg_4_ ( .D(n1609), .CK(CLK), .Q(node[4]) );
  DFFQX1 t12_reg_6_ ( .D(n1631), .CK(CLK), .Q(t12[6]) );
  DFFQX1 c22_reg_7_ ( .D(n1656), .CK(CLK), .Q(c22[7]) );
  DFFQX1 c12_reg_7_ ( .D(n1672), .CK(CLK), .Q(c12[7]) );
  DFFQX1 t21_reg_6_ ( .D(n1639), .CK(CLK), .Q(t21[6]) );
  DFFQX1 t22_reg_7_ ( .D(n1622), .CK(CLK), .Q(t22[7]) );
  DFFQX1 c12_reg_6_ ( .D(n1673), .CK(CLK), .Q(c12[6]) );
  DFFQX1 t11_reg_7_ ( .D(n1614), .CK(CLK), .Q(t11[7]) );
  DFFQX1 t22_reg_6_ ( .D(n1623), .CK(CLK), .Q(t22[6]) );
  DFFQX1 t12_reg_3_ ( .D(n1634), .CK(CLK), .Q(t12[3]) );
  DFFQX1 c12_reg_5_ ( .D(n1674), .CK(CLK), .Q(c12[5]) );
  DFFQX1 c12_reg_3_ ( .D(n1676), .CK(CLK), .Q(c12[3]) );
  DFFQX1 t12_reg_2_ ( .D(n1635), .CK(CLK), .Q(t12[2]) );
  DFFQX1 t21_reg_2_ ( .D(n1643), .CK(CLK), .Q(t21[2]) );
  DFFQX1 c12_reg_0_ ( .D(n1679), .CK(CLK), .Q(c12[0]) );
  DFFQX1 c21_reg_0_ ( .D(n1671), .CK(CLK), .Q(c21[0]) );
  DFFQX1 t12_reg_1_ ( .D(n1636), .CK(CLK), .Q(t12[1]) );
  DFFQX1 t21_reg_5_ ( .D(n1640), .CK(CLK), .Q(t21[5]) );
  DFFQX1 t22_reg_5_ ( .D(n1624), .CK(CLK), .Q(t22[5]) );
  DFFQX1 t22_reg_3_ ( .D(n1626), .CK(CLK), .Q(t22[3]) );
  DFFQX1 t21_reg_3_ ( .D(n1642), .CK(CLK), .Q(t21[3]) );
  DFFQX1 t11_reg_3_ ( .D(n1618), .CK(CLK), .Q(t11[3]) );
  DFFQX1 c22_reg_6_ ( .D(n1657), .CK(CLK), .Q(c22[6]) );
  DFFQX1 t12_reg_5_ ( .D(n1632), .CK(CLK), .Q(t12[5]) );
  DFFQX1 t11_reg_5_ ( .D(n1616), .CK(CLK), .Q(t11[5]) );
  DFFQX1 max12_reg_0_ ( .D(n1597), .CK(CLK), .Q(N1310) );
  DFFQX1 c11_reg_6_ ( .D(n1647), .CK(CLK), .Q(c11[6]) );
  DFFHQX8 out_reg_8_ ( .D(n1501), .CK(CLK), .Q(out[8]) );
  DFFHQX8 out_reg_2_ ( .D(n1507), .CK(CLK), .Q(out[2]) );
  DFFHQX8 out_reg_3_ ( .D(n1506), .CK(CLK), .Q(out[3]) );
  DFFHQX8 out_reg_4_ ( .D(n1505), .CK(CLK), .Q(out[4]) );
  DFFHQX8 out_reg_5_ ( .D(n1504), .CK(CLK), .Q(out[5]) );
  DFFHQX8 out_reg_6_ ( .D(n1503), .CK(CLK), .Q(out[6]) );
  DFFHQX8 out_reg_7_ ( .D(n1502), .CK(CLK), .Q(out[7]) );
  EDFFX1 out_reg_1_ ( .D(n3074), .E(n8330), .CK(CLK), .QN(n1894) );
  EDFFX1 out_reg_0_ ( .D(n3073), .E(n8330), .CK(CLK), .QN(n1892) );
  DFFTRX1 mode_reg_5_ ( .D(N154), .RN(n3075), .CK(CLK), .Q(mode[5]), .QN(n383)
         );
  DFFTRX1 mode_reg_2_ ( .D(N151), .RN(n3075), .CK(CLK), .Q(mode[2]), .QN(n388)
         );
  DFFTRX1 mode_reg_1_ ( .D(N150), .RN(n3075), .CK(CLK), .Q(mode[1]), .QN(n390)
         );
  DFFTRX1 mode_reg_7_ ( .D(N156), .RN(n3075), .CK(CLK), .Q(mode[7]), .QN(n2316) );
  DFFXL start_reg_0_ ( .D(N182), .CK(CLK), .Q(n2996), .QN(n398) );
  DFFXL a7_reg_8_ ( .D(n1517), .CK(CLK), .QN(n745) );
  DFFXL a7_reg_7_ ( .D(n1518), .CK(CLK), .Q(n2964), .QN(n746) );
  DFFXL a7_reg_6_ ( .D(n1519), .CK(CLK), .Q(n2962), .QN(n747) );
  DFFXL a7_reg_2_ ( .D(n1523), .CK(CLK), .Q(n2954), .QN(n751) );
  DFFXL a7_reg_0_ ( .D(n1525), .CK(CLK), .Q(n2948), .QN(n753) );
  DFFXL a5_reg_7_ ( .D(n1536), .CK(CLK), .Q(n2927), .QN(n763) );
  DFFXL a5_reg_6_ ( .D(n1537), .CK(CLK), .Q(n2925), .QN(n764) );
  DFFXL a5_reg_5_ ( .D(n1538), .CK(CLK), .Q(n2923), .QN(n765) );
  DFFXL a5_reg_4_ ( .D(n1539), .CK(CLK), .Q(n2921), .QN(n766) );
  DFFXL a5_reg_3_ ( .D(n1540), .CK(CLK), .Q(n2919), .QN(n767) );
  DFFXL a5_reg_2_ ( .D(n1541), .CK(CLK), .Q(n2917), .QN(n768) );
  DFFXL a5_reg_1_ ( .D(n1542), .CK(CLK), .Q(n2915), .QN(n769) );
  DFFXL a5_reg_0_ ( .D(n1543), .CK(CLK), .Q(n2911), .QN(n770) );
  DFFXL a4_reg_7_ ( .D(n1545), .CK(CLK), .Q(n2909), .QN(n754) );
  DFFXL a4_reg_6_ ( .D(n1546), .CK(CLK), .Q(n2907), .QN(n755) );
  DFFXL a4_reg_5_ ( .D(n1547), .CK(CLK), .Q(n2905), .QN(n756) );
  DFFXL a4_reg_4_ ( .D(n1548), .CK(CLK), .Q(n2903), .QN(n757) );
  DFFXL a4_reg_3_ ( .D(n1549), .CK(CLK), .Q(n2901), .QN(n758) );
  DFFXL a4_reg_2_ ( .D(n1550), .CK(CLK), .Q(n2899), .QN(n759) );
  DFFXL a4_reg_1_ ( .D(n1551), .CK(CLK), .Q(n2897), .QN(n760) );
  DFFXL a3_reg_7_ ( .D(n1554), .CK(CLK), .Q(n2891), .QN(n735) );
  DFFXL a3_reg_6_ ( .D(n1555), .CK(CLK), .Q(n2889), .QN(n736) );
  DFFXL a3_reg_5_ ( .D(n1556), .CK(CLK), .Q(n2887), .QN(n737) );
  DFFXL a3_reg_4_ ( .D(n1557), .CK(CLK), .Q(n2885), .QN(n738) );
  DFFXL a3_reg_3_ ( .D(n1558), .CK(CLK), .Q(n2883), .QN(n739) );
  DFFXL a3_reg_2_ ( .D(n1559), .CK(CLK), .Q(n2881), .QN(n740) );
  DFFXL a3_reg_1_ ( .D(n1560), .CK(CLK), .Q(n2879), .QN(n741) );
  DFFXL a3_reg_0_ ( .D(n1561), .CK(CLK), .Q(n2875), .QN(n742) );
  DFFXL a6_reg_7_ ( .D(n1527), .CK(CLK), .Q(n2945), .QN(n772) );
  DFFXL a6_reg_6_ ( .D(n1528), .CK(CLK), .Q(n2943), .QN(n773) );
  DFFXL a6_reg_5_ ( .D(n1529), .CK(CLK), .Q(n2941), .QN(n774) );
  DFFXL a6_reg_4_ ( .D(n1530), .CK(CLK), .Q(n2939), .QN(n775) );
  DFFXL a6_reg_3_ ( .D(n1531), .CK(CLK), .Q(n2937), .QN(n776) );
  DFFXL a6_reg_2_ ( .D(n1532), .CK(CLK), .Q(n2935), .QN(n777) );
  DFFXL a6_reg_1_ ( .D(n1533), .CK(CLK), .Q(n2933), .QN(n778) );
  DFFXL a6_reg_0_ ( .D(n1534), .CK(CLK), .Q(n2929), .QN(n779) );
  DFFXL a4_reg_0_ ( .D(n1552), .CK(CLK), .Q(n2893), .QN(n761) );
  DFFXL a1_reg_8_ ( .D(n1508), .CK(CLK), .QN(n780) );
  DFFXL a1_reg_7_ ( .D(n1509), .CK(CLK), .QN(n781) );
  DFFXL a1_reg_6_ ( .D(n1510), .CK(CLK), .QN(n782) );
  DFFXL a1_reg_5_ ( .D(n1511), .CK(CLK), .QN(n783) );
  DFFXL a1_reg_4_ ( .D(n1512), .CK(CLK), .QN(n784) );
  DFFXL a1_reg_3_ ( .D(n1513), .CK(CLK), .QN(n785) );
  DFFXL a1_reg_2_ ( .D(n1514), .CK(CLK), .QN(n786) );
  DFFXL a7_reg_5_ ( .D(n1520), .CK(CLK), .Q(n2960), .QN(n748) );
  DFFXL a7_reg_4_ ( .D(n1521), .CK(CLK), .Q(n2958), .QN(n749) );
  DFFXL a7_reg_3_ ( .D(n1522), .CK(CLK), .Q(n2956), .QN(n750) );
  DFFXL a7_reg_1_ ( .D(n1524), .CK(CLK), .Q(n2952), .QN(n752) );
  DFFQX1 t11_reg_4_ ( .D(n1617), .CK(CLK), .Q(t11[4]) );
  EDFFXL m65_reg_6_ ( .D(n3077), .E(n1445), .CK(CLK), .QN(n415) );
  EDFFXL m65_reg_5_ ( .D(n3078), .E(n1445), .CK(CLK), .QN(n416) );
  EDFFXL m65_reg_4_ ( .D(n3079), .E(n1445), .CK(CLK), .QN(n417) );
  EDFFXL m65_reg_3_ ( .D(n3080), .E(n1445), .CK(CLK), .QN(n418) );
  EDFFXL m65_reg_2_ ( .D(n3081), .E(n1445), .CK(CLK), .QN(n419) );
  EDFFXL m65_reg_1_ ( .D(n3082), .E(n1445), .CK(CLK), .QN(n420) );
  EDFFXL m63_reg_6_ ( .D(n3077), .E(n1450), .CK(CLK), .Q(n2466), .QN(n400) );
  EDFFXL m63_reg_5_ ( .D(n3078), .E(n1450), .CK(CLK), .Q(n2453), .QN(n401) );
  EDFFXL m63_reg_4_ ( .D(n3079), .E(n1450), .CK(CLK), .Q(n2440), .QN(n402) );
  EDFFXL m63_reg_3_ ( .D(n3080), .E(n1450), .CK(CLK), .Q(n2427), .QN(n403) );
  EDFFXL m63_reg_2_ ( .D(n3081), .E(n1450), .CK(CLK), .Q(n2414), .QN(n404) );
  EDFFXL m63_reg_1_ ( .D(n3082), .E(n1450), .CK(CLK), .Q(n2401), .QN(n405) );
  EDFFXL m62_reg_6_ ( .D(n3077), .E(n1452), .CK(CLK), .QN(n423) );
  EDFFXL m62_reg_5_ ( .D(n3078), .E(n1452), .CK(CLK), .QN(n424) );
  EDFFXL m62_reg_4_ ( .D(n3079), .E(n1452), .CK(CLK), .QN(n425) );
  EDFFXL m62_reg_3_ ( .D(n3080), .E(n1452), .CK(CLK), .QN(n426) );
  EDFFXL m62_reg_2_ ( .D(n3081), .E(n1452), .CK(CLK), .QN(n427) );
  EDFFXL m62_reg_1_ ( .D(n3082), .E(n1452), .CK(CLK), .QN(n428) );
  EDFFXL m62_reg_0_ ( .D(n3083), .E(n1452), .CK(CLK), .QN(n429) );
  EDFFXL m56_reg_6_ ( .D(n3077), .E(n1456), .CK(CLK), .QN(n674) );
  EDFFXL m56_reg_5_ ( .D(n3078), .E(n1456), .CK(CLK), .QN(n675) );
  EDFFXL m56_reg_4_ ( .D(n3079), .E(n1456), .CK(CLK), .QN(n676) );
  EDFFXL m56_reg_3_ ( .D(n3080), .E(n1456), .CK(CLK), .QN(n677) );
  EDFFXL m56_reg_2_ ( .D(n3081), .E(n1456), .CK(CLK), .QN(n678) );
  EDFFXL m56_reg_1_ ( .D(n3082), .E(n1456), .CK(CLK), .QN(n679) );
  EDFFXL m56_reg_0_ ( .D(n3083), .E(n1456), .CK(CLK), .QN(n680) );
  EDFFXL m13_reg_6_ ( .D(n3077), .E(n1490), .CK(CLK), .QN(n458) );
  EDFFXL m13_reg_5_ ( .D(n3078), .E(n1490), .CK(CLK), .QN(n459) );
  EDFFXL m13_reg_4_ ( .D(n3079), .E(n1490), .CK(CLK), .QN(n460) );
  EDFFXL m13_reg_3_ ( .D(n3080), .E(n1490), .CK(CLK), .QN(n461) );
  EDFFXL m13_reg_2_ ( .D(n3081), .E(n1490), .CK(CLK), .QN(n462) );
  EDFFXL m13_reg_1_ ( .D(n3082), .E(n1490), .CK(CLK), .QN(n463) );
  EDFFXL m66_reg_4_ ( .D(n3079), .E(n1443), .CK(CLK), .QN(n432) );
  EDFFXL m66_reg_2_ ( .D(n3081), .E(n1443), .CK(CLK), .QN(n434) );
  EDFFXL m61_reg_4_ ( .D(n3079), .E(n1454), .CK(CLK), .QN(n683) );
  EDFFXL m61_reg_2_ ( .D(n3081), .E(n1454), .CK(CLK), .QN(n685) );
  EDFFXL m65_reg_0_ ( .D(n3083), .E(n1445), .CK(CLK), .QN(n421) );
  EDFFXL m63_reg_0_ ( .D(n3083), .E(n1450), .CK(CLK), .Q(n2386), .QN(n406) );
  EDFFXL m13_reg_0_ ( .D(n3083), .E(n1490), .CK(CLK), .QN(n464) );
  EDFFXL m66_reg_6_ ( .D(n3077), .E(n1443), .CK(CLK), .QN(n430) );
  EDFFXL m66_reg_3_ ( .D(n3080), .E(n1443), .CK(CLK), .QN(n433) );
  EDFFXL m66_reg_1_ ( .D(n3082), .E(n1443), .CK(CLK), .QN(n435) );
  EDFFXL m66_reg_0_ ( .D(n3083), .E(n1443), .CK(CLK), .QN(n436) );
  EDFFXL m61_reg_6_ ( .D(n3077), .E(n1454), .CK(CLK), .QN(n681) );
  EDFFXL m61_reg_3_ ( .D(n3080), .E(n1454), .CK(CLK), .QN(n684) );
  EDFFXL m61_reg_1_ ( .D(n3082), .E(n1454), .CK(CLK), .QN(n686) );
  EDFFXL m61_reg_0_ ( .D(n3083), .E(n1454), .CK(CLK), .QN(n687) );
  EDFFXL m66_reg_5_ ( .D(n3078), .E(n1443), .CK(CLK), .QN(n431) );
  EDFFXL m61_reg_5_ ( .D(n3078), .E(n1454), .CK(CLK), .QN(n682) );
  DFFXL start_reg_1_ ( .D(N183), .CK(CLK), .Q(start_1_), .QN(n2997) );
  DFFTRX2 mode_reg_6_ ( .D(N155), .RN(n3075), .CK(CLK), .Q(n2785), .QN(n2317)
         );
  DFFTRX2 mode_reg_4_ ( .D(N153), .RN(n3075), .CK(CLK), .Q(mode[4]), .QN(n385)
         );
  DFFTRX2 mode_reg_0_ ( .D(N149), .RN(n3075), .CK(CLK), .Q(mode[0]), .QN(N1001) );
  DFFTRX2 mode_reg_3_ ( .D(N152), .RN(n3075), .CK(CLK), .Q(mode[3]), .QN(n386)
         );
  DFFQX1 max22_reg_7_ ( .D(n1574), .CK(CLK), .Q(max22[7]) );
  DFFQX1 max21_reg_0_ ( .D(n1589), .CK(CLK), .Q(N1329) );
  DFFQX1 max11_reg_0_ ( .D(n1605), .CK(CLK), .Q(N1291) );
  DFFQX1 max22_reg_0_ ( .D(n1581), .CK(CLK), .Q(N1348) );
  DFFQX1 t11_reg_6_ ( .D(n1615), .CK(CLK), .Q(t11[6]) );
  DFFQX1 t11_reg_2_ ( .D(n1619), .CK(CLK), .Q(t11[2]) );
  DFFQX1 t11_reg_1_ ( .D(n1620), .CK(CLK), .Q(t11[1]) );
  DFFQX1 t22_reg_4_ ( .D(n1625), .CK(CLK), .Q(t22[4]) );
  DFFQX1 t12_reg_7_ ( .D(n1630), .CK(CLK), .Q(t12[7]) );
  DFFQX1 c21_reg_6_ ( .D(n1665), .CK(CLK), .Q(c21[6]) );
  DFFQX1 s1_reg ( .D(n1573), .CK(CLK), .Q(s1) );
  DFFQX1 c22_reg_0_ ( .D(n1663), .CK(CLK), .Q(c22[0]) );
  DFFQX2 c11_reg_4_ ( .D(n1649), .CK(CLK), .Q(c11[4]) );
  DFFQX2 c11_reg_2_ ( .D(n1651), .CK(CLK), .Q(c11[2]) );
  DFFQX4 c22_reg_1_ ( .D(n1662), .CK(CLK), .Q(c22[1]) );
  DFFQX2 c22_reg_2_ ( .D(n1661), .CK(CLK), .Q(c22[2]) );
  DFFQX2 c12_reg_4_ ( .D(n1675), .CK(CLK), .Q(c12[4]) );
  DFFQX2 c22_reg_4_ ( .D(n1659), .CK(CLK), .Q(c22[4]) );
  DFFQX2 t22_reg_1_ ( .D(n1628), .CK(CLK), .Q(t22[1]) );
  DFFQX2 c21_reg_1_ ( .D(n1670), .CK(CLK), .Q(c21[1]) );
  DFFX2 t21_reg_0_ ( .D(n1645), .CK(CLK), .Q(n1898) );
  DFFQX2 t11_reg_0_ ( .D(n1621), .CK(CLK), .Q(t11[0]) );
  DFFQX2 c22_reg_3_ ( .D(n1660), .CK(CLK), .Q(c22[3]) );
  DFFQX2 t21_reg_4_ ( .D(n1641), .CK(CLK), .Q(t21[4]) );
  DFFQX2 t22_reg_2_ ( .D(n1627), .CK(CLK), .Q(t22[2]) );
  DFFQX2 c12_reg_2_ ( .D(n1677), .CK(CLK), .Q(c12[2]) );
  DFFQX2 c21_reg_3_ ( .D(n1668), .CK(CLK), .Q(c21[3]) );
  DFFQX2 c21_reg_2_ ( .D(n1669), .CK(CLK), .Q(c21[2]) );
  DFFQX2 t21_reg_1_ ( .D(n1644), .CK(CLK), .Q(t21[1]) );
  DFFQX2 t12_reg_4_ ( .D(n1633), .CK(CLK), .Q(t12[4]) );
  DFFQX2 c11_reg_0_ ( .D(n1653), .CK(CLK), .Q(c11[0]) );
  DFFQX2 t22_reg_0_ ( .D(n1629), .CK(CLK), .Q(t22[0]) );
  DFFQX2 c12_reg_1_ ( .D(n1678), .CK(CLK), .Q(c12[1]) );
  DFFQX2 t12_reg_0_ ( .D(n1637), .CK(CLK), .Q(t12[0]) );
  DFFQX2 c21_reg_4_ ( .D(n1667), .CK(CLK), .Q(c21[4]) );
  MXI2XL U1052 ( .A(N844), .B(N836), .S0(n1777), .Y(n2811) );
  MXI2XL U1053 ( .A(N845), .B(N837), .S0(n1777), .Y(n2812) );
  OA22X1 U1054 ( .A0(n2269), .A1(t22[3]), .B0(n2269), .B1(n2283), .Y(n2273) );
  NOR2BX1 U1055 ( .AN(t21[4]), .B(c21[4]), .Y(n2256) );
  CLKINVX1 U1056 ( .A(c12[1]), .Y(n2245) );
  OAI222X2 U1057 ( .A0(t12[5]), .A1(n2247), .B0(t12[5]), .B1(n2230), .C0(n2247), .C1(n2230), .Y(n2231) );
  INVX3 U1058 ( .A(n3003), .Y(n8330) );
  AOI21X1 U1059 ( .A0(t22[1]), .A1(n2282), .B0(t22[0]), .Y(n2270) );
  NOR2X1 U1060 ( .A(n2816), .B(n2148), .Y(n1929) );
  MXI2X2 U1061 ( .A(N868), .B(N860), .S0(N858), .Y(n2816) );
  INVX3 U1062 ( .A(n2815), .Y(N856) );
  NAND2BX1 U1063 ( .AN(t12[4]), .B(c12[4]), .Y(n2230) );
  AOI21X1 U1064 ( .A0(t21[1]), .A1(n2263), .B0(n1898), .Y(n2252) );
  NOR2BX4 U1065 ( .AN(t21[2]), .B(c21[2]), .Y(n2251) );
  NAND2BX1 U1066 ( .AN(t21[2]), .B(c21[2]), .Y(n2253) );
  NOR2BX2 U1067 ( .AN(t12[2]), .B(c12[2]), .Y(n2232) );
  NAND2BX1 U1068 ( .AN(t12[2]), .B(c12[2]), .Y(n2234) );
  NOR2BX2 U1069 ( .AN(t22[2]), .B(c22[2]), .Y(n2269) );
  NAND2BX1 U1070 ( .AN(t22[2]), .B(c22[2]), .Y(n2271) );
  INVX1 U1071 ( .A(c22[3]), .Y(n2283) );
  AOI2BB2X1 U1072 ( .B0(n2270), .B1(c22[0]), .A0N(t22[1]), .A1N(n2282), .Y(
        n2272) );
  CLKINVX8 U1073 ( .A(n2826), .Y(N904) );
  MXI2X4 U1074 ( .A(N896), .B(N888), .S0(N885), .Y(n2826) );
  MXI2X4 U1075 ( .A(N842), .B(N834), .S0(n1777), .Y(n2809) );
  NAND2BX2 U1076 ( .AN(t22[4]), .B(c22[4]), .Y(n2267) );
  NOR2BX1 U1077 ( .AN(t22[4]), .B(c22[4]), .Y(n2274) );
  INVX4 U1078 ( .A(n2808), .Y(N849) );
  OR2XL U1079 ( .A(n2808), .B(n2148), .Y(n1931) );
  MXI2X4 U1080 ( .A(N841), .B(N833), .S0(n1777), .Y(n2808) );
  MXI2X2 U1081 ( .A(N924), .B(N916), .S0(n2088), .Y(n2835) );
  CLKINVX1 U1082 ( .A(c22[1]), .Y(n2282) );
  OAI221X2 U1083 ( .A0(c12[6]), .A1(n2244), .B0(n2240), .B1(n2239), .C0(n2238), 
        .Y(n2241) );
  OAI22X2 U1084 ( .A0(n2236), .A1(n2235), .B0(n2234), .B1(n2246), .Y(n2239) );
  OAI22X1 U1085 ( .A0(t12[3]), .A1(n2246), .B0(t12[3]), .B1(n2234), .Y(n2240)
         );
  NOR2BX4 U1086 ( .AN(t11[2]), .B(c11[2]), .Y(n2213) );
  NAND2BX1 U1087 ( .AN(t11[2]), .B(c11[2]), .Y(n2215) );
  NOR2BX1 U1088 ( .AN(t11[4]), .B(c11[4]), .Y(n2218) );
  NAND2BX4 U1089 ( .AN(t11[4]), .B(c11[4]), .Y(n2211) );
  OAI222X1 U1090 ( .A0(N994), .A1(n2297), .B0(n2311), .B1(n2297), .C0(N994), 
        .C1(n2311), .Y(n2298) );
  OAI222X4 U1091 ( .A0(N963), .A1(n2306), .B0(N963), .B1(n2296), .C0(n2306), 
        .C1(n2296), .Y(n2297) );
  CLKINVX1 U1092 ( .A(n2824), .Y(N883) );
  CLKINVX1 U1093 ( .A(n2821), .Y(N880) );
  CLKINVX1 U1094 ( .A(n2812), .Y(N853) );
  NAND3X2 U1095 ( .A(n1960), .B(n1961), .C(n1962), .Y(n2287) );
  CLKINVX1 U1096 ( .A(t12[6]), .Y(n2244) );
  OR2X2 U1097 ( .A(n1918), .B(n1919), .Y(n2258) );
  OAI22X1 U1098 ( .A0(n2273), .A1(n2272), .B0(n2271), .B1(n2283), .Y(n2276) );
  CLKINVX1 U1099 ( .A(t22[6]), .Y(n2281) );
  MXI2X1 U1100 ( .A(N902), .B(N894), .S0(N885), .Y(n2832) );
  CLKINVX1 U1101 ( .A(n2822), .Y(N881) );
  CLKINVX1 U1102 ( .A(n2811), .Y(N852) );
  CLKINVX1 U1103 ( .A(n2820), .Y(N879) );
  CLKINVX1 U1104 ( .A(n2825), .Y(N903) );
  CLKINVX1 U1105 ( .A(c11[1]), .Y(n2226) );
  NAND2BX1 U1106 ( .AN(t21[4]), .B(c21[4]), .Y(n2249) );
  NAND3X1 U1107 ( .A(n1908), .B(n1909), .C(n1910), .Y(n2212) );
  CLKINVX1 U1108 ( .A(N997), .Y(n1903) );
  NOR2X1 U1109 ( .A(n2287), .B(n2312), .Y(n1958) );
  NOR2X1 U1110 ( .A(N997), .B(n2287), .Y(n1957) );
  OAI21XL U1111 ( .A0(n2300), .A1(n2299), .B0(n2298), .Y(n2302) );
  OR2X1 U1112 ( .A(n1933), .B(n1934), .Y(n2220) );
  OR2X4 U1113 ( .A(n2259), .B(n2258), .Y(n1921) );
  NOR2X1 U1114 ( .A(c21[6]), .B(n2250), .Y(n1926) );
  NAND3X1 U1115 ( .A(n1922), .B(n1923), .C(n2275), .Y(n2278) );
  OR3X2 U1116 ( .A(n1943), .B(n1944), .C(n1945), .Y(n2279) );
  NAND2X1 U1117 ( .A(n2304), .B(n2303), .Y(N999) );
  NAND2X1 U1118 ( .A(n2302), .B(n1950), .Y(n2303) );
  OR3X2 U1119 ( .A(n1957), .B(n1958), .C(n1959), .Y(n2304) );
  AOI21X1 U1120 ( .A0(n1903), .A1(N967), .B0(n1904), .Y(n1950) );
  NAND2X4 U1121 ( .A(N999), .B(n2682), .Y(n2807) );
  NAND2X1 U1122 ( .A(N914), .B(n2088), .Y(n1941) );
  NAND2X1 U1123 ( .A(N922), .B(n1939), .Y(n1940) );
  MXI2X1 U1124 ( .A(N929), .B(N921), .S0(n2088), .Y(n2840) );
  OR4X1 U1125 ( .A(n2672), .B(n2673), .C(n2674), .D(n2675), .Y(n1897) );
  NAND2X1 U1126 ( .A(N928), .B(n1914), .Y(n1915) );
  BUFX2 U1127 ( .A(n2178), .Y(n2177) );
  OR2X1 U1128 ( .A(n2825), .B(n2148), .Y(n1924) );
  NAND3X1 U1129 ( .A(n1912), .B(n1913), .C(n2170), .Y(n1574) );
  OR2X1 U1130 ( .A(n2149), .B(n2210), .Y(n1913) );
  OR2X1 U1131 ( .A(n2840), .B(n2148), .Y(n1912) );
  NAND2X1 U1132 ( .A(n1901), .B(n1902), .Y(n1573) );
  NAND3X1 U1133 ( .A(n1899), .B(n1900), .C(n2173), .Y(n1582) );
  OR2X1 U1134 ( .A(n2832), .B(n2148), .Y(n1899) );
  BUFX12 U1135 ( .A(n1949), .Y(n2149) );
  NAND2X6 U1136 ( .A(n2170), .B(n2807), .Y(n1949) );
  INVX3 U1137 ( .A(n2348), .Y(n2365) );
  INVX3 U1138 ( .A(n2177), .Y(n2170) );
  NAND2X1 U1139 ( .A(n2780), .B(n2778), .Y(n1683) );
  NAND3X1 U1140 ( .A(n2784), .B(n2785), .C(n2351), .Y(n1684) );
  NAND2XL U1141 ( .A(n2789), .B(n2780), .Y(n1685) );
  NAND2X1 U1142 ( .A(n2782), .B(n2780), .Y(n1686) );
  NAND2X1 U1143 ( .A(n2354), .B(n2782), .Y(n1687) );
  NAND2X1 U1144 ( .A(n2359), .B(n2782), .Y(n1688) );
  OR2X1 U1145 ( .A(n2177), .B(n2323), .Y(n1697) );
  NAND2X1 U1146 ( .A(n2782), .B(n2351), .Y(n1698) );
  NAND2X1 U1147 ( .A(n2778), .B(n2779), .Y(n1699) );
  NAND2XL U1148 ( .A(n2789), .B(n2779), .Y(n1700) );
  NAND3X1 U1149 ( .A(n2784), .B(n2785), .C(n2783), .Y(n1701) );
  OA21XL U1150 ( .A0(n2790), .A1(n3055), .B0(n2174), .Y(n1734) );
  NAND2X1 U1151 ( .A(n2789), .B(n2359), .Y(n1735) );
  NAND2XL U1152 ( .A(n2789), .B(n2357), .Y(n1736) );
  NAND2X1 U1153 ( .A(n2782), .B(n2783), .Y(n1737) );
  NAND2X1 U1154 ( .A(n2789), .B(n2781), .Y(n1738) );
  NAND2X1 U1155 ( .A(n2782), .B(n2779), .Y(n1739) );
  NAND2X1 U1156 ( .A(n2357), .B(n2782), .Y(n1740) );
  NAND2X1 U1157 ( .A(n2781), .B(n2778), .Y(n1741) );
  OA21XL U1158 ( .A0(n2791), .A1(n3055), .B0(n2173), .Y(n1774) );
  OA21XL U1159 ( .A0(n2360), .A1(n2790), .B0(n2173), .Y(n1775) );
  OA21XL U1160 ( .A0(n2360), .A1(n2791), .B0(n2173), .Y(n1776) );
  CLKINVX1 U1161 ( .A(c21[1]), .Y(n2263) );
  CLKINVX1 U1162 ( .A(n1942), .Y(n2833) );
  NAND2X1 U1163 ( .A(n1940), .B(n1941), .Y(n1942) );
  CLKINVX1 U1164 ( .A(c21[5]), .Y(n2265) );
  NAND2X1 U1165 ( .A(n2682), .B(n2149), .Y(n1952) );
  OAI21X4 U1166 ( .A0(t11[7]), .A1(n2229), .B0(n2224), .Y(n1777) );
  NAND2X4 U1167 ( .A(n1935), .B(n2243), .Y(N858) );
  CLKINVX1 U1168 ( .A(n1917), .Y(n2839) );
  CLKINVX1 U1169 ( .A(N1310), .Y(n2817) );
  CLKINVX1 U1170 ( .A(max22[1]), .Y(n2204) );
  NAND2X1 U1171 ( .A(sub_516_S2_carry[7]), .B(n2187), .Y(n1778) );
  NAND2X1 U1172 ( .A(sub_518_S2_carry[7]), .B(n2194), .Y(n1779) );
  NAND2X1 U1173 ( .A(sub_520_S2_carry[7]), .B(n2202), .Y(n1780) );
  NAND2X1 U1174 ( .A(sub_522_S2_carry[7]), .B(n2210), .Y(n1781) );
  CLKINVX1 U1175 ( .A(N1348), .Y(n2203) );
  NOR3X1 U1176 ( .A(mode[4]), .B(mode[5]), .C(mode[3]), .Y(n2784) );
  OAI21X2 U1177 ( .A0(n2367), .A1(n3058), .B0(n2174), .Y(n1458) );
  AND2X2 U1178 ( .A(in[0]), .B(n2365), .Y(n3083) );
  AND2X2 U1179 ( .A(in[1]), .B(n2365), .Y(n3082) );
  AND2X2 U1180 ( .A(in[2]), .B(n2365), .Y(n3081) );
  AND2X2 U1181 ( .A(in[3]), .B(n2365), .Y(n3080) );
  AND2X2 U1182 ( .A(in[4]), .B(n2365), .Y(n3079) );
  AND2X2 U1183 ( .A(in[5]), .B(n2365), .Y(n3078) );
  AND2X2 U1184 ( .A(in[6]), .B(n2365), .Y(n3077) );
  NOR3XL U1185 ( .A(mode[3]), .B(n383), .C(mode[4]), .Y(n3062) );
  INVX3 U1186 ( .A(n1776), .Y(n1838) );
  INVX3 U1187 ( .A(n1775), .Y(n1839) );
  INVX3 U1188 ( .A(n1774), .Y(n1840) );
  INVX3 U1189 ( .A(n1734), .Y(n1841) );
  OAI21X2 U1190 ( .A0(n3058), .A1(n2790), .B0(n2174), .Y(n1448) );
  OAI21X2 U1191 ( .A0(n3052), .A1(n3058), .B0(n2174), .Y(n1459) );
  OAI21X2 U1192 ( .A0(n2790), .A1(n3053), .B0(n2173), .Y(n1483) );
  OAI21X2 U1193 ( .A0(n3058), .A1(n2793), .B0(n2174), .Y(n1456) );
  OAI21X2 U1194 ( .A0(n2795), .A1(n3053), .B0(n2173), .Y(n1485) );
  NAND2X2 U1195 ( .A(n3061), .B(mode[0]), .Y(n2797) );
  OAI21X2 U1196 ( .A0(n3058), .A1(n2795), .B0(n2174), .Y(n1452) );
  OAI21X2 U1197 ( .A0(n2793), .A1(n3053), .B0(n2173), .Y(n1487) );
  OAI21X2 U1198 ( .A0(n3058), .A1(n2797), .B0(n2174), .Y(n1445) );
  OAI21X2 U1199 ( .A0(n3052), .A1(n3053), .B0(n2173), .Y(n1489) );
  NOR2X2 U1200 ( .A(n2091), .B(s4), .Y(n2930) );
  OAI21X2 U1201 ( .A0(n2797), .A1(n3053), .B0(n2173), .Y(n1481) );
  OAI21X2 U1202 ( .A0(n2795), .A1(n3055), .B0(n2174), .Y(n1475) );
  OAI21X2 U1203 ( .A0(n3052), .A1(n3057), .B0(n2171), .Y(n1469) );
  NOR2X2 U1204 ( .A(n2177), .B(n2089), .Y(n2684) );
  NOR2X2 U1205 ( .A(n2091), .B(s3), .Y(n2912) );
  OAI21X2 U1206 ( .A0(n2360), .A1(n2797), .B0(n2172), .Y(n1490) );
  NAND2X1 U1207 ( .A(n2365), .B(n2350), .Y(n2360) );
  OAI21X2 U1208 ( .A0(n3058), .A1(n2791), .B0(n2174), .Y(n1450) );
  OAI21X2 U1209 ( .A0(n2793), .A1(n3055), .B0(n2173), .Y(n1477) );
  OAI21X2 U1210 ( .A0(n3057), .A1(n2790), .B0(n2174), .Y(n1463) );
  NAND2X2 U1211 ( .A(n2170), .B(n3063), .Y(n1443) );
  INVX3 U1212 ( .A(n1970), .Y(n2338) );
  NOR2X2 U1213 ( .A(n2091), .B(s2), .Y(n2894) );
  MXI2X2 U1214 ( .A(n2177), .B(N999), .S0(n2682), .Y(n2805) );
  OA21X2 U1215 ( .A0(n2354), .A1(n2179), .B0(n1911), .Y(n2353) );
  OAI21X2 U1216 ( .A0(n2367), .A1(n3053), .B0(n2172), .Y(n1488) );
  OAI21X2 U1217 ( .A0(n2797), .A1(n3055), .B0(n2173), .Y(n1471) );
  OAI21X2 U1218 ( .A0(n3057), .A1(n2795), .B0(n2174), .Y(n1465) );
  NAND2BX2 U1219 ( .AN(n2994), .B(n2323), .Y(n2873) );
  INVX3 U1220 ( .A(n3032), .Y(n2339) );
  INVX6 U1221 ( .A(n1892), .Y(out[0]) );
  NOR2X2 U1222 ( .A(mode[0]), .B(n2803), .Y(n2351) );
  NOR2X2 U1223 ( .A(n2091), .B(s1), .Y(n2876) );
  OA21X2 U1224 ( .A0(n2359), .A1(n2177), .B0(n1911), .Y(n2358) );
  OAI21X2 U1225 ( .A0(n2791), .A1(n3053), .B0(n2172), .Y(n1484) );
  OAI21X2 U1226 ( .A0(n2794), .A1(n3055), .B0(n2173), .Y(n1476) );
  OAI21X2 U1227 ( .A0(n3057), .A1(n2793), .B0(n2174), .Y(n1467) );
  NAND2X2 U1228 ( .A(n2348), .B(n2349), .Y(n3075) );
  INVX3 U1229 ( .A(n3031), .Y(n2340) );
  INVX3 U1230 ( .A(node[4]), .Y(n2325) );
  INVX6 U1231 ( .A(n1894), .Y(out[1]) );
  OAI211XL U1232 ( .A0(n3021), .A1(n2999), .B0(n3022), .C0(n3023), .Y(n1503)
         );
  OAI211XL U1233 ( .A0(n3016), .A1(n2999), .B0(n3017), .C0(n3018), .Y(n1504)
         );
  OAI211XL U1234 ( .A0(n3011), .A1(n2999), .B0(n3012), .C0(n3013), .Y(n1505)
         );
  OAI211XL U1235 ( .A0(n3006), .A1(n2999), .B0(n3007), .C0(n3008), .Y(n1506)
         );
  OAI211XL U1236 ( .A0(n2998), .A1(n2999), .B0(n3000), .C0(n3001), .Y(n1507)
         );
  OAI211XL U1237 ( .A0(n3033), .A1(n2999), .B0(n3034), .C0(n3035), .Y(n1501)
         );
  NOR3X2 U1238 ( .A(node[6]), .B(node[7]), .C(node[5]), .Y(n2333) );
  NOR2X2 U1239 ( .A(n2965), .B(n2091), .Y(n2949) );
  OA21X2 U1240 ( .A0(n2994), .A1(n2972), .B0(n2986), .Y(n2991) );
  NAND3XL U1241 ( .A(n2995), .B(n2352), .C(n2170), .Y(n2972) );
  OA21X2 U1242 ( .A0(n2357), .A1(n2176), .B0(n2355), .Y(n2356) );
  NAND2XL U1243 ( .A(n2170), .B(n2360), .Y(n2355) );
  OA21X2 U1244 ( .A0(in_valid), .A1(n2177), .B0(n2366), .Y(n2364) );
  OAI21X2 U1245 ( .A0(n2794), .A1(n3053), .B0(n2172), .Y(n1486) );
  OAI21X2 U1246 ( .A0(n3052), .A1(n3055), .B0(n2173), .Y(n1479) );
  OAI21X2 U1247 ( .A0(n3057), .A1(n2797), .B0(n2174), .Y(n1461) );
  AOI31X1 U1248 ( .A0(n2682), .A1(n1897), .A2(n2316), .B0(n2176), .Y(n1896) );
  INVX3 U1249 ( .A(n2831), .Y(N909) );
  OR2XL U1250 ( .A(n2149), .B(n2202), .Y(n1900) );
  OR2X1 U1251 ( .A(n2149), .B(n2841), .Y(n1901) );
  OR2XL U1252 ( .A(n1777), .B(n2148), .Y(n1902) );
  OA22X2 U1253 ( .A0(n2301), .A1(n2307), .B0(n2301), .B1(N966), .Y(n1904) );
  NOR2X1 U1254 ( .A(c11[6]), .B(n2212), .Y(n1905) );
  NOR2X1 U1255 ( .A(n2225), .B(n2212), .Y(n1906) );
  NOR2X1 U1256 ( .A(c11[6]), .B(n2225), .Y(n1907) );
  OR3X2 U1257 ( .A(n1905), .B(n1906), .C(n1907), .Y(n2223) );
  OR2X1 U1258 ( .A(t11[5]), .B(n2228), .Y(n1908) );
  OR2X2 U1259 ( .A(t11[5]), .B(n2211), .Y(n1909) );
  OR2X2 U1260 ( .A(n2228), .B(n2211), .Y(n1910) );
  CLKINVX1 U1261 ( .A(t11[6]), .Y(n2225) );
  AO22X4 U1262 ( .A0(n2229), .A1(t11[7]), .B0(n2223), .B1(n2222), .Y(n2224) );
  INVX4 U1263 ( .A(c11[5]), .Y(n2228) );
  NAND2XL U1264 ( .A(n2170), .B(n2360), .Y(n1911) );
  CLKINVX2 U1265 ( .A(n2807), .Y(n2806) );
  OR2X4 U1266 ( .A(n2286), .B(n2307), .Y(n1962) );
  OR2X4 U1267 ( .A(N966), .B(n2286), .Y(n1961) );
  NAND2BX1 U1268 ( .AN(N965), .B(N995), .Y(n2286) );
  NAND2X1 U1269 ( .A(N920), .B(n2088), .Y(n1916) );
  NAND2X1 U1270 ( .A(n1915), .B(n1916), .Y(n1917) );
  INVXL U1271 ( .A(n2088), .Y(n1914) );
  BUFX20 U1272 ( .A(N912), .Y(n2088) );
  NOR2X1 U1273 ( .A(n2255), .B(n2254), .Y(n1918) );
  NOR2X1 U1274 ( .A(n2253), .B(n2264), .Y(n1919) );
  OR2X1 U1275 ( .A(c21[6]), .B(n2262), .Y(n1920) );
  NAND3X4 U1276 ( .A(n1920), .B(n1921), .C(n2257), .Y(n2260) );
  AOI2BB2XL U1277 ( .B0(n2252), .B1(c21[0]), .A0N(t21[1]), .A1N(n2263), .Y(
        n2254) );
  CLKINVX1 U1278 ( .A(c21[3]), .Y(n2264) );
  AOI22X4 U1279 ( .A0(n2266), .A1(t21[7]), .B0(n2261), .B1(n2260), .Y(n1954)
         );
  OR2X4 U1280 ( .A(n2277), .B(n2276), .Y(n1923) );
  NOR2X1 U1281 ( .A(n2262), .B(n2250), .Y(n1927) );
  OR3X2 U1282 ( .A(n1926), .B(n1927), .C(n1928), .Y(n2261) );
  MX2XL U1283 ( .A(c11[4]), .B(n2160), .S0(n2364), .Y(n1649) );
  INVX1 U1284 ( .A(n2819), .Y(N878) );
  OAI221X1 U1285 ( .A0(c11[6]), .A1(n2225), .B0(n2221), .B1(n2220), .C0(n2219), 
        .Y(n2222) );
  NAND3X1 U1286 ( .A(n1924), .B(n1925), .C(n2174), .Y(n1589) );
  OR2XL U1287 ( .A(n2149), .B(n2195), .Y(n1925) );
  AOI2BB2X2 U1288 ( .B0(n2214), .B1(c11[0]), .A0N(t11[1]), .A1N(n2226), .Y(
        n2216) );
  INVX1 U1289 ( .A(t21[6]), .Y(n2262) );
  NOR2X1 U1290 ( .A(c21[6]), .B(n2262), .Y(n1928) );
  INVX4 U1291 ( .A(n1963), .Y(n2250) );
  OR2XL U1292 ( .A(c22[6]), .B(n2281), .Y(n1922) );
  AO22X4 U1293 ( .A0(n2285), .A1(t22[7]), .B0(n2279), .B1(n2278), .Y(n2280) );
  BUFX12 U1294 ( .A(n1952), .Y(n2148) );
  NOR2XL U1295 ( .A(n2215), .B(n2227), .Y(n1934) );
  NOR2X4 U1296 ( .A(n2217), .B(n2216), .Y(n1933) );
  AOI21X4 U1297 ( .A0(t11[1]), .A1(n2226), .B0(t11[0]), .Y(n2214) );
  NAND3X1 U1298 ( .A(n1931), .B(n1932), .C(n2172), .Y(n1605) );
  CLKINVX1 U1299 ( .A(c22[7]), .Y(n2285) );
  OR2X1 U1300 ( .A(t12[7]), .B(n2248), .Y(n1935) );
  MXI2X2 U1301 ( .A(N895), .B(N887), .S0(N885), .Y(n2825) );
  CLKINVX3 U1302 ( .A(N962), .Y(n2310) );
  INVX3 U1303 ( .A(n2176), .Y(n2172) );
  OR3X2 U1304 ( .A(n1929), .B(n1930), .C(n2179), .Y(n1597) );
  OAI21X4 U1305 ( .A0(t22[7]), .A1(n2285), .B0(n2280), .Y(N912) );
  INVX1 U1306 ( .A(c12[7]), .Y(n2248) );
  INVX4 U1307 ( .A(c11[3]), .Y(n2227) );
  NOR2XL U1308 ( .A(n2149), .B(n2817), .Y(n1930) );
  OR2X1 U1309 ( .A(n2149), .B(n2180), .Y(n1932) );
  MX2XL U1310 ( .A(c11[2]), .B(n2164), .S0(n2364), .Y(n1651) );
  NOR2BX1 U1311 ( .AN(t12[4]), .B(c12[4]), .Y(n2237) );
  OA22X2 U1312 ( .A0(n2232), .A1(t12[3]), .B0(n2232), .B1(n2246), .Y(n2236) );
  INVX3 U1313 ( .A(n2088), .Y(n1939) );
  INVX1 U1314 ( .A(n2351), .Y(n3052) );
  OR2XL U1315 ( .A(t22[5]), .B(n2284), .Y(n1946) );
  OR2XL U1316 ( .A(c12[6]), .B(n2244), .Y(n1938) );
  INVX8 U1317 ( .A(n1953), .Y(N885) );
  MXI2XL U1318 ( .A(N927), .B(N919), .S0(n2088), .Y(n2838) );
  MXI2XL U1319 ( .A(N925), .B(N917), .S0(n2088), .Y(n2836) );
  MXI2XL U1320 ( .A(N926), .B(N918), .S0(n2088), .Y(n2837) );
  NOR2X1 U1321 ( .A(c22[6]), .B(n2268), .Y(n1943) );
  NOR2X1 U1322 ( .A(n2281), .B(n2268), .Y(n1944) );
  OR2X1 U1323 ( .A(t22[5]), .B(n2267), .Y(n1947) );
  OR2X1 U1324 ( .A(n2284), .B(n2267), .Y(n1948) );
  NAND3X2 U1325 ( .A(n1946), .B(n1947), .C(n1948), .Y(n2268) );
  OR2X1 U1326 ( .A(c12[6]), .B(n2231), .Y(n1936) );
  OR2X1 U1327 ( .A(n2244), .B(n2231), .Y(n1937) );
  NAND3X1 U1328 ( .A(n1936), .B(n1937), .C(n1938), .Y(n2242) );
  AO22X4 U1329 ( .A0(n2248), .A1(t12[7]), .B0(n2242), .B1(n2241), .Y(n2243) );
  NOR2BX1 U1330 ( .AN(N965), .B(N995), .Y(n2301) );
  CLKINVX1 U1331 ( .A(n3041), .Y(n2328) );
  OR2X1 U1332 ( .A(N966), .B(n2307), .Y(n1960) );
  NOR2X1 U1333 ( .A(n2310), .B(N992), .Y(n2294) );
  INVX3 U1334 ( .A(n2814), .Y(N855) );
  AND4X1 U1335 ( .A(n3043), .B(N1073), .C(N1075), .D(N1074), .Y(n1680) );
  AND2X2 U1336 ( .A(n2796), .B(mode[3]), .Y(n2782) );
  AND2XL U1337 ( .A(n2778), .B(n2351), .Y(n2384) );
  NAND3XL U1338 ( .A(n2850), .B(n2325), .C(n2990), .Y(n2870) );
  INVXL U1339 ( .A(n2333), .Y(n2345) );
  NAND3XL U1340 ( .A(n2850), .B(n2325), .C(n2872), .Y(n2858) );
  INVX3 U1341 ( .A(n2249), .Y(n1965) );
  INVX3 U1342 ( .A(t21[5]), .Y(n1964) );
  OAI22XL U1343 ( .A0(n2256), .A1(n2265), .B0(t21[5]), .B1(n2256), .Y(n2257)
         );
  AOI21X1 U1344 ( .A0(t12[1]), .A1(n2245), .B0(t12[0]), .Y(n2233) );
  OA22X2 U1345 ( .A0(n2251), .A1(t21[3]), .B0(n2251), .B1(n2264), .Y(n2255) );
  OA22X2 U1346 ( .A0(n2213), .A1(t11[3]), .B0(n2213), .B1(n2227), .Y(n2217) );
  CLKINVX1 U1347 ( .A(finish), .Y(n1955) );
  AOI32XL U1348 ( .A0(n2985), .A1(n2344), .A2(n2333), .B0(n2974), .B1(a1[1]), 
        .Y(n2984) );
  AND2X2 U1349 ( .A(n2796), .B(n386), .Y(n2778) );
  INVX3 U1350 ( .A(c22[5]), .Y(n2284) );
  NOR2X1 U1351 ( .A(c22[6]), .B(n2281), .Y(n1945) );
  INVX1 U1352 ( .A(N964), .Y(n2311) );
  INVXL U1353 ( .A(n2290), .Y(n2309) );
  INVX3 U1354 ( .A(n2823), .Y(N882) );
  INVX3 U1355 ( .A(n2813), .Y(N854) );
  INVX3 U1356 ( .A(n2810), .Y(N851) );
  AND2XL U1357 ( .A(n2995), .B(n2328), .Y(n2986) );
  CLKBUFX2 U1358 ( .A(n2179), .Y(n2175) );
  NOR2X1 U1359 ( .A(n2671), .B(n1896), .Y(n1951) );
  CLKINVX1 U1360 ( .A(N996), .Y(n2307) );
  INVX3 U1361 ( .A(n2816), .Y(N876) );
  OAI211XL U1362 ( .A0(n2850), .A1(n2857), .B0(n2872), .C0(n2325), .Y(n2871)
         );
  AOI2BB1XL U1363 ( .A0N(n3067), .A1N(n3041), .B0(n3064), .Y(N182) );
  AOI2BB1X4 U1364 ( .A0N(t21[7]), .A1N(n2266), .B0(n1954), .Y(n1953) );
  INVX3 U1365 ( .A(c12[5]), .Y(n2247) );
  INVX3 U1366 ( .A(c12[3]), .Y(n2246) );
  NAND2X8 U1367 ( .A(n1955), .B(n1956), .Y(n1969) );
  CLKINVX20 U1368 ( .A(RESET), .Y(n1956) );
  NOR3X2 U1369 ( .A(n398), .B(start_1_), .C(n2176), .Y(n2682) );
  NAND2XL U1370 ( .A(out[8]), .B(n3003), .Y(n3034) );
  NAND2XL U1371 ( .A(out[2]), .B(n3003), .Y(n3000) );
  NAND2XL U1372 ( .A(out[3]), .B(n3003), .Y(n3007) );
  NAND2XL U1373 ( .A(out[4]), .B(n3003), .Y(n3012) );
  NAND2XL U1374 ( .A(out[5]), .B(n3003), .Y(n3017) );
  NAND2XL U1375 ( .A(out[6]), .B(n3003), .Y(n3022) );
  NAND2XL U1376 ( .A(out[7]), .B(n3003), .Y(n3027) );
  MXI2XL U1377 ( .A(n2318), .B(n2319), .S0(n2320), .Y(n3072) );
  OAI32XL U1378 ( .A0(n2324), .A1(node[0]), .A2(n2325), .B0(node[2]), .B1(
        n2326), .Y(n2322) );
  MXI2XL U1379 ( .A(n2845), .B(n2846), .S0(n2320), .Y(n1569) );
  AO22XL U1380 ( .A0(t21[5]), .A1(n2095), .B0(n2097), .B1(n2441), .Y(n1640) );
  AO22XL U1381 ( .A0(t12[5]), .A1(n2095), .B0(n2096), .B1(n2539), .Y(n1632) );
  AO22XL U1382 ( .A0(t22[5]), .A1(n2095), .B0(n2096), .B1(n2635), .Y(n1624) );
  AO22XL U1383 ( .A0(t21[3]), .A1(n2095), .B0(n2097), .B1(n2415), .Y(n1642) );
  AO22XL U1384 ( .A0(t12[3]), .A1(n2095), .B0(n2097), .B1(n2515), .Y(n1634) );
  AO22XL U1385 ( .A0(t22[3]), .A1(n2095), .B0(n2096), .B1(n2611), .Y(n1626) );
  AO22XL U1386 ( .A0(n1898), .A1(n2095), .B0(n2097), .B1(n2368), .Y(n1645) );
  AO22XL U1387 ( .A0(t12[0]), .A1(n2095), .B0(n2097), .B1(n2479), .Y(n1637) );
  AO22XL U1388 ( .A0(t22[0]), .A1(n2095), .B0(n2096), .B1(n2575), .Y(n1629) );
  AO22XL U1389 ( .A0(t21[1]), .A1(n2095), .B0(n2097), .B1(n2389), .Y(n1644) );
  AO22XL U1390 ( .A0(t12[1]), .A1(n2095), .B0(n2097), .B1(n2491), .Y(n1636) );
  AO22XL U1391 ( .A0(t22[1]), .A1(n2095), .B0(n2096), .B1(n2587), .Y(n1628) );
  AO22XL U1392 ( .A0(t21[7]), .A1(n2095), .B0(n2097), .B1(n2467), .Y(n1638) );
  AO22XL U1393 ( .A0(t12[7]), .A1(n2095), .B0(n2096), .B1(n2563), .Y(n1630) );
  AO22XL U1394 ( .A0(t22[7]), .A1(n2095), .B0(n2096), .B1(n2659), .Y(n1622) );
  AO22XL U1395 ( .A0(t21[2]), .A1(n2095), .B0(n2097), .B1(n2402), .Y(n1643) );
  AO22XL U1396 ( .A0(t12[2]), .A1(n2095), .B0(n2097), .B1(n2503), .Y(n1635) );
  AO22XL U1397 ( .A0(t12[4]), .A1(n1896), .B0(n2096), .B1(n2527), .Y(n1633) );
  AO22XL U1398 ( .A0(t22[2]), .A1(n1896), .B0(n2096), .B1(n2599), .Y(n1627) );
  AO22XL U1399 ( .A0(t22[4]), .A1(n2095), .B0(n2096), .B1(n2623), .Y(n1625) );
  AO22XL U1400 ( .A0(t21[4]), .A1(n2095), .B0(n2097), .B1(n2428), .Y(n1641) );
  AO22XL U1401 ( .A0(t21[6]), .A1(n2095), .B0(n2097), .B1(n2454), .Y(n1639) );
  AO22XL U1402 ( .A0(t12[6]), .A1(n1896), .B0(n2096), .B1(n2551), .Y(n1631) );
  AO22XL U1403 ( .A0(t22[6]), .A1(n2095), .B0(n2096), .B1(n2647), .Y(n1623) );
  MX2XL U1404 ( .A(c21[0]), .B(n2168), .S0(n2356), .Y(n1671) );
  MX2XL U1405 ( .A(c21[1]), .B(n2166), .S0(n2356), .Y(n1670) );
  MX2XL U1406 ( .A(c21[2]), .B(n2164), .S0(n2356), .Y(n1669) );
  MX2XL U1407 ( .A(c21[3]), .B(n2162), .S0(n2356), .Y(n1668) );
  MX2XL U1408 ( .A(c21[4]), .B(n2160), .S0(n2356), .Y(n1667) );
  MX2XL U1409 ( .A(c21[6]), .B(n2156), .S0(n2356), .Y(n1665) );
  MX2XL U1410 ( .A(c21[7]), .B(n2154), .S0(n2356), .Y(n1664) );
  MX2XL U1411 ( .A(c12[0]), .B(n2168), .S0(n2353), .Y(n1679) );
  MX2XL U1412 ( .A(c12[1]), .B(n2166), .S0(n2353), .Y(n1678) );
  MX2XL U1413 ( .A(c12[2]), .B(n2164), .S0(n2353), .Y(n1677) );
  MX2XL U1414 ( .A(c12[3]), .B(n2162), .S0(n2353), .Y(n1676) );
  MX2XL U1415 ( .A(c12[4]), .B(n2160), .S0(n2353), .Y(n1675) );
  MX2XL U1416 ( .A(c12[5]), .B(n2158), .S0(n2353), .Y(n1674) );
  MX2XL U1417 ( .A(c12[6]), .B(n2156), .S0(n2353), .Y(n1673) );
  MX2XL U1418 ( .A(c12[7]), .B(n2154), .S0(n2353), .Y(n1672) );
  MX2XL U1419 ( .A(c22[0]), .B(n2168), .S0(n2358), .Y(n1663) );
  MX2XL U1420 ( .A(c22[1]), .B(n2166), .S0(n2358), .Y(n1662) );
  MX2XL U1421 ( .A(c22[2]), .B(n2164), .S0(n2358), .Y(n1661) );
  MX2XL U1422 ( .A(c22[3]), .B(n2162), .S0(n2358), .Y(n1660) );
  MX2XL U1423 ( .A(c22[4]), .B(n2160), .S0(n2358), .Y(n1659) );
  MX2XL U1424 ( .A(c22[5]), .B(n2158), .S0(n2358), .Y(n1658) );
  MX2XL U1425 ( .A(c22[6]), .B(n2156), .S0(n2358), .Y(n1657) );
  MX2XL U1426 ( .A(c22[7]), .B(n2154), .S0(n2358), .Y(n1656) );
  MX2XL U1427 ( .A(n2331), .B(n2332), .S0(n2333), .Y(n2330) );
  XNOR2XL U1428 ( .A(N1291), .B(N1329), .Y(n2969) );
  INVXL U1429 ( .A(max21[1]), .Y(n2196) );
  INVXL U1430 ( .A(max11[1]), .Y(n2181) );
  INVXL U1431 ( .A(max12[1]), .Y(n2188) );
  XNOR2XL U1432 ( .A(max11[1]), .B(n2971), .Y(n2966) );
  XNOR3XL U1433 ( .A(n2204), .B(max21[1]), .C(max12[1]), .Y(n2967) );
  INVXL U1434 ( .A(max12[2]), .Y(n2189) );
  INVXL U1435 ( .A(max22[2]), .Y(n2205) );
  INVXL U1436 ( .A(max11[2]), .Y(n2182) );
  INVXL U1437 ( .A(max21[2]), .Y(n2197) );
  INVXL U1438 ( .A(N1291), .Y(n2180) );
  INVXL U1439 ( .A(N1329), .Y(n2195) );
  INVXL U1440 ( .A(max12[3]), .Y(n2190) );
  INVXL U1441 ( .A(max22[3]), .Y(n2206) );
  INVXL U1442 ( .A(max21[3]), .Y(n2198) );
  NOR2XL U1443 ( .A(N1348), .B(N1310), .Y(n2970) );
  NAND2XL U1444 ( .A(N1329), .B(N1291), .Y(n2971) );
  NOR2X1 U1445 ( .A(N997), .B(n2312), .Y(n1959) );
  AOI222X4 U1446 ( .A0(n1964), .A1(c21[5]), .B0(n1964), .B1(n1965), .C0(c21[5]), .C1(n1965), .Y(n1963) );
  CLKBUFX3 U1447 ( .A(n2385), .Y(n2143) );
  CLKINVX1 U1448 ( .A(N959), .Y(n2308) );
  INVX3 U1449 ( .A(n2153), .Y(n2150) );
  INVX3 U1450 ( .A(n2153), .Y(n2151) );
  CLKINVX1 U1451 ( .A(n2153), .Y(n2152) );
  CLKBUFX3 U1452 ( .A(n2109), .Y(n2108) );
  CLKBUFX3 U1453 ( .A(n2118), .Y(n2119) );
  CLKBUFX3 U1454 ( .A(n2112), .Y(n2113) );
  CLKBUFX3 U1455 ( .A(n2104), .Y(n2105) );
  CLKBUFX3 U1456 ( .A(n2114), .Y(n2115) );
  CLKBUFX3 U1457 ( .A(n2385), .Y(n2142) );
  CLKBUFX3 U1458 ( .A(n1697), .Y(n2153) );
  CLKINVX1 U1459 ( .A(N967), .Y(n2312) );
  CLKBUFX3 U1460 ( .A(n1951), .Y(n2097) );
  CLKBUFX3 U1461 ( .A(n1951), .Y(n2096) );
  AND2X2 U1462 ( .A(n2873), .B(n2153), .Y(n2320) );
  INVX3 U1463 ( .A(n2176), .Y(n2173) );
  CLKBUFX3 U1464 ( .A(n3076), .Y(n2155) );
  INVX3 U1465 ( .A(n2175), .Y(n2174) );
  CLKBUFX3 U1466 ( .A(n1686), .Y(n2118) );
  CLKBUFX3 U1467 ( .A(n1687), .Y(n2104) );
  CLKBUFX3 U1468 ( .A(n1688), .Y(n2114) );
  CLKBUFX3 U1469 ( .A(n2111), .Y(n2110) );
  CLKBUFX3 U1470 ( .A(n1739), .Y(n2111) );
  CLKBUFX3 U1471 ( .A(n2384), .Y(n2141) );
  CLKBUFX3 U1472 ( .A(n2127), .Y(n2126) );
  CLKBUFX3 U1473 ( .A(n2123), .Y(n2122) );
  CLKBUFX3 U1474 ( .A(n1683), .Y(n2101) );
  CLKBUFX3 U1475 ( .A(n1685), .Y(n2133) );
  CLKBUFX3 U1476 ( .A(n1741), .Y(n2099) );
  CLKBUFX3 U1477 ( .A(n2103), .Y(n2102) );
  CLKBUFX3 U1478 ( .A(n2135), .Y(n2134) );
  CLKBUFX3 U1479 ( .A(n2383), .Y(n2139) );
  CLKBUFX3 U1480 ( .A(n2125), .Y(n2124) );
  CLKBUFX3 U1481 ( .A(n1698), .Y(n2109) );
  CLKBUFX3 U1482 ( .A(n1740), .Y(n2112) );
  INVX3 U1483 ( .A(n2175), .Y(n2171) );
  CLKBUFX3 U1484 ( .A(n2146), .Y(n2147) );
  CLKBUFX3 U1485 ( .A(n2106), .Y(n2107) );
  CLKBUFX3 U1486 ( .A(n2117), .Y(n2116) );
  CLKBUFX3 U1487 ( .A(n2144), .Y(n2145) );
  CLKBUFX3 U1488 ( .A(n2136), .Y(n2137) );
  CLKBUFX3 U1489 ( .A(n2141), .Y(n2140) );
  CLKBUFX3 U1490 ( .A(n2133), .Y(n2132) );
  CLKBUFX3 U1491 ( .A(n2101), .Y(n2100) );
  CLKBUFX3 U1492 ( .A(n1741), .Y(n2098) );
  INVX3 U1493 ( .A(n2087), .Y(n1466) );
  CLKBUFX3 U1494 ( .A(n2179), .Y(n2176) );
  CLKBUFX3 U1495 ( .A(n2329), .Y(n2091) );
  CLKBUFX3 U1496 ( .A(n1896), .Y(n2095) );
  OAI21X2 U1497 ( .A0(n3057), .A1(n2367), .B0(n2174), .Y(n1468) );
  CLKBUFX3 U1498 ( .A(n3083), .Y(n2168) );
  CLKBUFX3 U1499 ( .A(n3082), .Y(n2166) );
  CLKBUFX3 U1500 ( .A(n3081), .Y(n2164) );
  CLKBUFX3 U1501 ( .A(n3080), .Y(n2162) );
  CLKBUFX3 U1502 ( .A(n3079), .Y(n2160) );
  CLKBUFX3 U1503 ( .A(n3078), .Y(n2158) );
  CLKBUFX3 U1504 ( .A(n3077), .Y(n2156) );
  CLKBUFX3 U1505 ( .A(n3083), .Y(n2169) );
  CLKBUFX3 U1506 ( .A(n3082), .Y(n2167) );
  CLKBUFX3 U1507 ( .A(n3081), .Y(n2165) );
  CLKBUFX3 U1508 ( .A(n3080), .Y(n2163) );
  CLKBUFX3 U1509 ( .A(n3079), .Y(n2161) );
  CLKBUFX3 U1510 ( .A(n3078), .Y(n2159) );
  CLKBUFX3 U1511 ( .A(n3077), .Y(n2157) );
  CLKBUFX3 U1512 ( .A(n3076), .Y(n2154) );
  CLKBUFX3 U1513 ( .A(n1737), .Y(n2106) );
  CLKBUFX3 U1514 ( .A(n2387), .Y(n2144) );
  CLKBUFX3 U1515 ( .A(n2382), .Y(n2136) );
  CLKBUFX3 U1516 ( .A(n2388), .Y(n2146) );
  CLKBUFX3 U1517 ( .A(n1738), .Y(n2135) );
  CLKBUFX3 U1518 ( .A(n1700), .Y(n2130) );
  CLKBUFX3 U1519 ( .A(n1735), .Y(n2123) );
  CLKBUFX3 U1520 ( .A(n2380), .Y(n2125) );
  CLKBUFX3 U1521 ( .A(n1736), .Y(n2127) );
  CLKBUFX3 U1522 ( .A(n2381), .Y(n2129) );
  CLKBUFX3 U1523 ( .A(n1699), .Y(n2103) );
  CLKINVX1 U1524 ( .A(N993), .Y(n2306) );
  CLKINVX1 U1525 ( .A(N991), .Y(n2305) );
  CLKBUFX3 U1526 ( .A(n2121), .Y(n2120) );
  CLKBUFX3 U1527 ( .A(n1684), .Y(n2121) );
  CLKBUFX3 U1528 ( .A(n2383), .Y(n2138) );
  CLKBUFX3 U1529 ( .A(n2129), .Y(n2128) );
  CLKBUFX3 U1530 ( .A(n1700), .Y(n2131) );
  CLKBUFX3 U1531 ( .A(n1701), .Y(n2117) );
  NOR4X2 U1532 ( .A(n2997), .B(n2996), .C(n2175), .D(n2094), .Y(n2323) );
  CLKBUFX3 U1533 ( .A(n1969), .Y(n2178) );
  CLKBUFX3 U1534 ( .A(n1969), .Y(n2179) );
  NOR2X2 U1535 ( .A(n2844), .B(n2091), .Y(n2931) );
  NOR2X2 U1536 ( .A(n2841), .B(n2091), .Y(n2877) );
  NOR2X2 U1537 ( .A(n2842), .B(n2091), .Y(n2895) );
  NOR2X2 U1538 ( .A(n2843), .B(n2091), .Y(n2913) );
  CLKBUFX3 U1539 ( .A(n2950), .Y(n2090) );
  NOR2BX1 U1540 ( .AN(n2965), .B(n2091), .Y(n2950) );
  AND2X2 U1541 ( .A(n2789), .B(n2354), .Y(n1966) );
  CLKINVX1 U1542 ( .A(n1966), .Y(n2380) );
  AND2X2 U1543 ( .A(n2789), .B(n2783), .Y(n1967) );
  CLKINVX1 U1544 ( .A(n1967), .Y(n2381) );
  NAND3X2 U1545 ( .A(N1075), .B(n3048), .C(N1073), .Y(n2337) );
  CLKINVX1 U1546 ( .A(c11[7]), .Y(n2229) );
  CLKINVX1 U1547 ( .A(c21[7]), .Y(n2266) );
  CLKBUFX3 U1548 ( .A(n2683), .Y(n2089) );
  CLKINVX1 U1549 ( .A(n2798), .Y(n2683) );
  CLKBUFX6 U1550 ( .A(n3113), .Y(out_valid) );
  NAND3X2 U1551 ( .A(N1075), .B(n3048), .C(outmode[0]), .Y(n2341) );
  CLKBUFX3 U1552 ( .A(n2334), .Y(n2092) );
  CLKBUFX3 U1553 ( .A(n3113), .Y(n2094) );
  AND3X2 U1554 ( .A(N1075), .B(N1074), .C(outmode[0]), .Y(n1970) );
  CLKINVX1 U1555 ( .A(max11[3]), .Y(n2183) );
  CLKINVX1 U1556 ( .A(max12[4]), .Y(n2191) );
  CLKINVX1 U1557 ( .A(max12[5]), .Y(n2192) );
  CLKINVX1 U1558 ( .A(max12[6]), .Y(n2193) );
  CLKINVX1 U1559 ( .A(max22[4]), .Y(n2207) );
  CLKINVX1 U1560 ( .A(max22[5]), .Y(n2208) );
  CLKINVX1 U1561 ( .A(max22[6]), .Y(n2209) );
  CLKINVX1 U1562 ( .A(max11[4]), .Y(n2184) );
  CLKINVX1 U1563 ( .A(max11[5]), .Y(n2185) );
  CLKINVX1 U1564 ( .A(max11[6]), .Y(n2186) );
  CLKINVX1 U1565 ( .A(max21[4]), .Y(n2199) );
  CLKINVX1 U1566 ( .A(max21[5]), .Y(n2200) );
  CLKINVX1 U1567 ( .A(max21[6]), .Y(n2201) );
  CLKINVX1 U1568 ( .A(max12[7]), .Y(n2194) );
  CLKINVX1 U1569 ( .A(max22[7]), .Y(n2210) );
  CLKINVX1 U1570 ( .A(max11[7]), .Y(n2187) );
  CLKINVX1 U1571 ( .A(max21[7]), .Y(n2202) );
  OAI21X2 U1572 ( .A0(n3058), .A1(n2794), .B0(n2171), .Y(n1454) );
  NAND3X2 U1573 ( .A(n2365), .B(n2801), .C(n3062), .Y(n3058) );
  NAND4X2 U1574 ( .A(n3056), .B(n2365), .C(n386), .D(mode[4]), .Y(n3055) );
  OAI21X2 U1575 ( .A0(n2367), .A1(n3055), .B0(n2173), .Y(n1478) );
  NAND2X2 U1576 ( .A(n3054), .B(mode[4]), .Y(n3057) );
  AND3X2 U1577 ( .A(n3056), .B(n2365), .C(mode[3]), .Y(n3054) );
  NAND2X2 U1578 ( .A(n3054), .B(n385), .Y(n3053) );
  OAI21X2 U1579 ( .A0(n3057), .A1(n2791), .B0(n2174), .Y(n1464) );
  AOI2BB1XL U1580 ( .A0N(n3057), .A1N(n2794), .B0(n2176), .Y(n2087) );
  INVXL U1581 ( .A(n2323), .Y(n2329) );
  AOI211X4 U1582 ( .A0(n3042), .A1(n3043), .B0(n1680), .C0(n2153), .Y(n3003)
         );
  MXI2XL U1583 ( .A(n2363), .B(n2362), .S0(n1458), .Y(n1654) );
  XOR2X1 U1584 ( .A(n2187), .B(sub_516_S2_carry[7]), .Y(N1298) );
  AND2X1 U1585 ( .A(sub_516_S2_carry[6]), .B(n2186), .Y(sub_516_S2_carry[7])
         );
  XOR2X1 U1586 ( .A(n2186), .B(sub_516_S2_carry[6]), .Y(N1297) );
  AND2X1 U1587 ( .A(sub_516_S2_carry[5]), .B(n2185), .Y(sub_516_S2_carry[6])
         );
  XOR2X1 U1588 ( .A(n2185), .B(sub_516_S2_carry[5]), .Y(N1296) );
  AND2X1 U1589 ( .A(sub_516_S2_carry[4]), .B(n2184), .Y(sub_516_S2_carry[5])
         );
  XOR2X1 U1590 ( .A(n2184), .B(sub_516_S2_carry[4]), .Y(N1295) );
  AND2X1 U1591 ( .A(sub_516_S2_carry[3]), .B(n2183), .Y(sub_516_S2_carry[4])
         );
  XOR2X1 U1592 ( .A(n2183), .B(sub_516_S2_carry[3]), .Y(N1294) );
  AND2X1 U1593 ( .A(sub_516_S2_carry[2]), .B(n2182), .Y(sub_516_S2_carry[3])
         );
  XOR2X1 U1594 ( .A(n2182), .B(sub_516_S2_carry[2]), .Y(N1293) );
  AND2X1 U1595 ( .A(n2180), .B(n2181), .Y(sub_516_S2_carry[2]) );
  XOR2X1 U1596 ( .A(n2181), .B(n2180), .Y(N1292) );
  XOR2X1 U1597 ( .A(n2194), .B(sub_518_S2_carry[7]), .Y(N1317) );
  AND2X1 U1598 ( .A(sub_518_S2_carry[6]), .B(n2193), .Y(sub_518_S2_carry[7])
         );
  XOR2X1 U1599 ( .A(n2193), .B(sub_518_S2_carry[6]), .Y(N1316) );
  AND2X1 U1600 ( .A(sub_518_S2_carry[5]), .B(n2192), .Y(sub_518_S2_carry[6])
         );
  XOR2X1 U1601 ( .A(n2192), .B(sub_518_S2_carry[5]), .Y(N1315) );
  AND2X1 U1602 ( .A(sub_518_S2_carry[4]), .B(n2191), .Y(sub_518_S2_carry[5])
         );
  XOR2X1 U1603 ( .A(n2191), .B(sub_518_S2_carry[4]), .Y(N1314) );
  AND2X1 U1604 ( .A(sub_518_S2_carry[3]), .B(n2190), .Y(sub_518_S2_carry[4])
         );
  XOR2X1 U1605 ( .A(n2190), .B(sub_518_S2_carry[3]), .Y(N1313) );
  AND2X1 U1606 ( .A(sub_518_S2_carry[2]), .B(n2189), .Y(sub_518_S2_carry[3])
         );
  XOR2X1 U1607 ( .A(n2189), .B(sub_518_S2_carry[2]), .Y(N1312) );
  AND2X1 U1608 ( .A(n2817), .B(n2188), .Y(sub_518_S2_carry[2]) );
  XOR2X1 U1609 ( .A(n2188), .B(n2817), .Y(N1311) );
  XOR2X1 U1610 ( .A(n2202), .B(sub_520_S2_carry[7]), .Y(N1336) );
  AND2X1 U1611 ( .A(sub_520_S2_carry[6]), .B(n2201), .Y(sub_520_S2_carry[7])
         );
  XOR2X1 U1612 ( .A(n2201), .B(sub_520_S2_carry[6]), .Y(N1335) );
  AND2X1 U1613 ( .A(sub_520_S2_carry[5]), .B(n2200), .Y(sub_520_S2_carry[6])
         );
  XOR2X1 U1614 ( .A(n2200), .B(sub_520_S2_carry[5]), .Y(N1334) );
  AND2X1 U1615 ( .A(sub_520_S2_carry[4]), .B(n2199), .Y(sub_520_S2_carry[5])
         );
  XOR2X1 U1616 ( .A(n2199), .B(sub_520_S2_carry[4]), .Y(N1333) );
  AND2X1 U1617 ( .A(sub_520_S2_carry[3]), .B(n2198), .Y(sub_520_S2_carry[4])
         );
  XOR2X1 U1618 ( .A(n2198), .B(sub_520_S2_carry[3]), .Y(N1332) );
  AND2X1 U1619 ( .A(sub_520_S2_carry[2]), .B(n2197), .Y(sub_520_S2_carry[3])
         );
  XOR2X1 U1620 ( .A(n2197), .B(sub_520_S2_carry[2]), .Y(N1331) );
  AND2X1 U1621 ( .A(n2195), .B(n2196), .Y(sub_520_S2_carry[2]) );
  XOR2X1 U1622 ( .A(n2196), .B(n2195), .Y(N1330) );
  XOR2X1 U1623 ( .A(n2210), .B(sub_522_S2_carry[7]), .Y(N1355) );
  AND2X1 U1624 ( .A(sub_522_S2_carry[6]), .B(n2209), .Y(sub_522_S2_carry[7])
         );
  XOR2X1 U1625 ( .A(n2209), .B(sub_522_S2_carry[6]), .Y(N1354) );
  AND2X1 U1626 ( .A(sub_522_S2_carry[5]), .B(n2208), .Y(sub_522_S2_carry[6])
         );
  XOR2X1 U1627 ( .A(n2208), .B(sub_522_S2_carry[5]), .Y(N1353) );
  AND2X1 U1628 ( .A(sub_522_S2_carry[4]), .B(n2207), .Y(sub_522_S2_carry[5])
         );
  XOR2X1 U1629 ( .A(n2207), .B(sub_522_S2_carry[4]), .Y(N1352) );
  AND2X1 U1630 ( .A(sub_522_S2_carry[3]), .B(n2206), .Y(sub_522_S2_carry[4])
         );
  XOR2X1 U1631 ( .A(n2206), .B(sub_522_S2_carry[3]), .Y(N1351) );
  AND2X1 U1632 ( .A(sub_522_S2_carry[2]), .B(n2205), .Y(sub_522_S2_carry[3])
         );
  XOR2X1 U1633 ( .A(n2205), .B(sub_522_S2_carry[2]), .Y(N1350) );
  AND2X1 U1634 ( .A(n2203), .B(n2204), .Y(sub_522_S2_carry[2]) );
  XOR2X1 U1635 ( .A(n2204), .B(n2203), .Y(N1349) );
  XNOR2X1 U1636 ( .A(mode[7]), .B(sub_404_carry_7_), .Y(N1008) );
  OR2X1 U1637 ( .A(n2785), .B(sub_404_carry_6_), .Y(sub_404_carry_7_) );
  XNOR2X1 U1638 ( .A(sub_404_carry_6_), .B(n2785), .Y(N1007) );
  AND2X1 U1639 ( .A(sub_404_carry_5_), .B(mode[5]), .Y(sub_404_carry_6_) );
  XOR2X1 U1640 ( .A(mode[5]), .B(sub_404_carry_5_), .Y(N1006) );
  OR2X1 U1641 ( .A(mode[4]), .B(sub_404_carry_4_), .Y(sub_404_carry_5_) );
  XNOR2X1 U1642 ( .A(sub_404_carry_4_), .B(mode[4]), .Y(N1005) );
  AND2X1 U1643 ( .A(sub_404_carry_3_), .B(mode[3]), .Y(sub_404_carry_4_) );
  XOR2X1 U1644 ( .A(mode[3]), .B(sub_404_carry_3_), .Y(N1004) );
  OR2X1 U1645 ( .A(mode[2]), .B(sub_404_carry_2_), .Y(sub_404_carry_3_) );
  XNOR2X1 U1646 ( .A(sub_404_carry_2_), .B(mode[2]), .Y(N1003) );
  OR2X1 U1647 ( .A(mode[1]), .B(mode[0]), .Y(sub_404_carry_2_) );
  XNOR2X1 U1648 ( .A(mode[0]), .B(mode[1]), .Y(N1002) );
  OAI22XL U1649 ( .A0(t11[3]), .A1(n2227), .B0(t11[3]), .B1(n2215), .Y(n2221)
         );
  OAI22XL U1650 ( .A0(n2218), .A1(n2228), .B0(t11[5]), .B1(n2218), .Y(n2219)
         );
  AOI2BB2X1 U1651 ( .B0(n2233), .B1(c12[0]), .A0N(t12[1]), .A1N(n2245), .Y(
        n2235) );
  OAI22XL U1652 ( .A0(n2237), .A1(n2247), .B0(t12[5]), .B1(n2237), .Y(n2238)
         );
  OAI22XL U1653 ( .A0(t21[3]), .A1(n2264), .B0(t21[3]), .B1(n2253), .Y(n2259)
         );
  OAI22XL U1654 ( .A0(t22[3]), .A1(n2283), .B0(t22[3]), .B1(n2271), .Y(n2277)
         );
  OAI22XL U1655 ( .A0(n2274), .A1(n2284), .B0(t22[5]), .B1(n2274), .Y(n2275)
         );
  NAND2BX1 U1656 ( .AN(N960), .B(N990), .Y(n2290) );
  AOI2BB1X1 U1657 ( .A0N(n2308), .A1N(N989), .B0(N958), .Y(n2288) );
  AO22X1 U1658 ( .A0(n2288), .A1(N988), .B0(N989), .B1(n2308), .Y(n2293) );
  NOR2BX1 U1659 ( .AN(N960), .B(N990), .Y(n2289) );
  OAI22XL U1660 ( .A0(n2289), .A1(n2305), .B0(N961), .B1(n2289), .Y(n2292) );
  OAI22XL U1661 ( .A0(N961), .A1(n2305), .B0(N961), .B1(n2290), .Y(n2291) );
  AOI221XL U1662 ( .A0(N991), .A1(n2309), .B0(n2293), .B1(n2292), .C0(n2291), 
        .Y(n2300) );
  OAI22XL U1663 ( .A0(n2294), .A1(n2306), .B0(N963), .B1(n2294), .Y(n2295) );
  OAI21XL U1664 ( .A0(N994), .A1(n2311), .B0(n2295), .Y(n2299) );
  NAND2X1 U1665 ( .A(N992), .B(n2310), .Y(n2296) );
  OAI21XL U1666 ( .A0(n2321), .A1(n2322), .B0(n2323), .Y(n2319) );
  CLKINVX1 U1667 ( .A(a2[0]), .Y(n2318) );
  OAI22XL U1668 ( .A0(n2327), .A1(n2328), .B0(n2091), .B1(n2330), .Y(n3073) );
  AOI211X1 U1669 ( .A0(n2092), .A1(a2[0]), .B0(n2335), .C0(n2336), .Y(n2327)
         );
  OAI22XL U1670 ( .A0(n779), .A1(n2337), .B0(n753), .B1(n2338), .Y(n2336) );
  OAI222XL U1671 ( .A0(n742), .A1(n2339), .B0(n761), .B1(n2340), .C0(n770), 
        .C1(n2341), .Y(n2335) );
  OAI22XL U1672 ( .A0(n2342), .A1(n2328), .B0(n2091), .B1(n2343), .Y(n3074) );
  MXI2X1 U1673 ( .A(n2344), .B(a1[1]), .S0(n2345), .Y(n2343) );
  AOI211X1 U1674 ( .A0(a2[1]), .A1(n2092), .B0(n2346), .C0(n2347), .Y(n2342)
         );
  OAI22XL U1675 ( .A0(n778), .A1(n2337), .B0(n752), .B1(n2338), .Y(n2347) );
  OAI222XL U1676 ( .A0(n741), .A1(n2339), .B0(n760), .B1(n2340), .C0(n769), 
        .C1(n2341), .Y(n2346) );
  OAI2BB1X1 U1677 ( .A0N(n2350), .A1N(n2351), .B0(n2170), .Y(n2349) );
  OAI31XL U1678 ( .A0(n2153), .A1(n1680), .A2(n2352), .B0(n2091), .Y(n1681) );
  CLKMX2X2 U1679 ( .A(c21[5]), .B(n2158), .S0(n2356), .Y(n1666) );
  MXI2X1 U1680 ( .A(n2361), .B(n2362), .S0(n1468), .Y(n1655) );
  CLKMX2X2 U1681 ( .A(c11[0]), .B(n2168), .S0(n2364), .Y(n1653) );
  CLKMX2X2 U1682 ( .A(c11[1]), .B(n2166), .S0(n2364), .Y(n1652) );
  CLKMX2X2 U1683 ( .A(c11[3]), .B(n2162), .S0(n2364), .Y(n1650) );
  CLKMX2X2 U1684 ( .A(c11[5]), .B(n2158), .S0(n2364), .Y(n1648) );
  CLKMX2X2 U1685 ( .A(c11[6]), .B(n2156), .S0(n2364), .Y(n1647) );
  CLKMX2X2 U1686 ( .A(c11[7]), .B(n2154), .S0(n2364), .Y(n1646) );
  OAI21XL U1687 ( .A0(n2367), .A1(n2360), .B0(n2365), .Y(n2366) );
  CLKINVX1 U1688 ( .A(n2362), .Y(n3076) );
  NAND2X1 U1689 ( .A(in[7]), .B(n2365), .Y(n2362) );
  NAND4X1 U1690 ( .A(n2369), .B(n2370), .C(n2371), .D(n2372), .Y(n2368) );
  NOR4X1 U1691 ( .A(n2373), .B(n2374), .C(n2375), .D(n2376), .Y(n2372) );
  OAI222XL U1692 ( .A0(n624), .A1(n2098), .B0(n616), .B1(n2100), .C0(n608), 
        .C1(n2102), .Y(n2376) );
  OAI222XL U1693 ( .A0(n656), .A1(n2105), .B0(n648), .B1(n2107), .C0(n640), 
        .C1(n2108), .Y(n2375) );
  OAI222XL U1694 ( .A0(n687), .A1(n2110), .B0(n664), .B1(n2113), .C0(n672), 
        .C1(n2115), .Y(n2374) );
  OAI222XL U1695 ( .A0(n421), .A1(n2116), .B0(n429), .B1(n2119), .C0(n414), 
        .C1(n2120), .Y(n2373) );
  NOR3X1 U1696 ( .A(n2377), .B(n2378), .C(n2379), .Y(n2371) );
  OAI22XL U1697 ( .A0(n520), .A1(n2122), .B0(n504), .B1(n2125), .Y(n2379) );
  OAI22XL U1698 ( .A0(n512), .A1(n2126), .B0(n496), .B1(n2128), .Y(n2378) );
  OAI222XL U1699 ( .A0(n528), .A1(n2131), .B0(n544), .B1(n2132), .C0(n552), 
        .C1(n2134), .Y(n2377) );
  AOI222XL U1700 ( .A0(n2137), .A1(n1702), .B0(n2138), .B1(n1742), .C0(n2140), 
        .C1(n1689), .Y(n2370) );
  AOI222XL U1701 ( .A0(n2143), .A1(n2386), .B0(n2145), .B1(n1718), .C0(n2147), 
        .C1(n1822), .Y(n2369) );
  NAND4X1 U1702 ( .A(n2390), .B(n2391), .C(n2392), .D(n2393), .Y(n2389) );
  NOR4X1 U1703 ( .A(n2394), .B(n2395), .C(n2396), .D(n2397), .Y(n2393) );
  OAI222XL U1704 ( .A0(n623), .A1(n2098), .B0(n615), .B1(n2101), .C0(n607), 
        .C1(n2103), .Y(n2397) );
  OAI222XL U1705 ( .A0(n655), .A1(n2104), .B0(n647), .B1(n2106), .C0(n639), 
        .C1(n2108), .Y(n2396) );
  OAI222XL U1706 ( .A0(n686), .A1(n2110), .B0(n663), .B1(n2112), .C0(n671), 
        .C1(n2114), .Y(n2395) );
  OAI222XL U1707 ( .A0(n420), .A1(n1701), .B0(n428), .B1(n2118), .C0(n413), 
        .C1(n2120), .Y(n2394) );
  NOR3X1 U1708 ( .A(n2398), .B(n2399), .C(n2400), .Y(n2392) );
  OAI22XL U1709 ( .A0(n519), .A1(n2122), .B0(n503), .B1(n2380), .Y(n2400) );
  OAI22XL U1710 ( .A0(n511), .A1(n2127), .B0(n495), .B1(n2128), .Y(n2399) );
  OAI222XL U1711 ( .A0(n527), .A1(n2130), .B0(n543), .B1(n2133), .C0(n551), 
        .C1(n2134), .Y(n2398) );
  AOI222XL U1712 ( .A0(n2136), .A1(n1703), .B0(n2138), .B1(n1743), .C0(n2141), 
        .C1(n1690), .Y(n2391) );
  AOI222XL U1713 ( .A0(n2143), .A1(n2401), .B0(n2144), .B1(n1719), .C0(n2146), 
        .C1(n1823), .Y(n2390) );
  NAND4X1 U1714 ( .A(n2403), .B(n2404), .C(n2405), .D(n2406), .Y(n2402) );
  NOR4X1 U1715 ( .A(n2407), .B(n2408), .C(n2409), .D(n2410), .Y(n2406) );
  OAI222XL U1716 ( .A0(n622), .A1(n2098), .B0(n614), .B1(n2101), .C0(n606), 
        .C1(n2103), .Y(n2410) );
  OAI222XL U1717 ( .A0(n654), .A1(n2104), .B0(n646), .B1(n2106), .C0(n638), 
        .C1(n2109), .Y(n2409) );
  OAI222XL U1718 ( .A0(n685), .A1(n2110), .B0(n662), .B1(n2112), .C0(n670), 
        .C1(n2114), .Y(n2408) );
  OAI222XL U1719 ( .A0(n419), .A1(n1701), .B0(n427), .B1(n2118), .C0(n412), 
        .C1(n2120), .Y(n2407) );
  NOR3X1 U1720 ( .A(n2411), .B(n2412), .C(n2413), .Y(n2405) );
  OAI22XL U1721 ( .A0(n518), .A1(n2123), .B0(n502), .B1(n2125), .Y(n2413) );
  OAI22XL U1722 ( .A0(n510), .A1(n2127), .B0(n494), .B1(n2128), .Y(n2412) );
  OAI222XL U1723 ( .A0(n526), .A1(n2131), .B0(n542), .B1(n2133), .C0(n550), 
        .C1(n2135), .Y(n2411) );
  AOI222XL U1724 ( .A0(n2136), .A1(n1704), .B0(n2138), .B1(n1744), .C0(n2140), 
        .C1(n1691), .Y(n2404) );
  AOI222XL U1725 ( .A0(n2143), .A1(n2414), .B0(n2144), .B1(n1720), .C0(n2146), 
        .C1(n1824), .Y(n2403) );
  NAND4X1 U1726 ( .A(n2416), .B(n2417), .C(n2418), .D(n2419), .Y(n2415) );
  NOR4X1 U1727 ( .A(n2420), .B(n2421), .C(n2422), .D(n2423), .Y(n2419) );
  OAI222XL U1728 ( .A0(n621), .A1(n2098), .B0(n613), .B1(n2100), .C0(n605), 
        .C1(n1699), .Y(n2423) );
  OAI222XL U1729 ( .A0(n653), .A1(n2104), .B0(n645), .B1(n2106), .C0(n637), 
        .C1(n2109), .Y(n2422) );
  OAI222XL U1730 ( .A0(n684), .A1(n2110), .B0(n661), .B1(n2112), .C0(n669), 
        .C1(n2114), .Y(n2421) );
  OAI222XL U1731 ( .A0(n418), .A1(n1701), .B0(n426), .B1(n2118), .C0(n411), 
        .C1(n2120), .Y(n2420) );
  NOR3X1 U1732 ( .A(n2424), .B(n2425), .C(n2426), .Y(n2418) );
  OAI22XL U1733 ( .A0(n517), .A1(n2123), .B0(n501), .B1(n2125), .Y(n2426) );
  OAI22XL U1734 ( .A0(n509), .A1(n2127), .B0(n493), .B1(n2128), .Y(n2425) );
  OAI222XL U1735 ( .A0(n525), .A1(n2131), .B0(n541), .B1(n2132), .C0(n549), 
        .C1(n2135), .Y(n2424) );
  AOI222XL U1736 ( .A0(n2136), .A1(n1705), .B0(n2138), .B1(n1745), .C0(n2140), 
        .C1(n1692), .Y(n2417) );
  AOI222XL U1737 ( .A0(n2143), .A1(n2427), .B0(n2144), .B1(n1721), .C0(n2146), 
        .C1(n1825), .Y(n2416) );
  NAND4X1 U1738 ( .A(n2429), .B(n2430), .C(n2431), .D(n2432), .Y(n2428) );
  NOR4X1 U1739 ( .A(n2433), .B(n2434), .C(n2435), .D(n2436), .Y(n2432) );
  OAI222XL U1740 ( .A0(n620), .A1(n2098), .B0(n612), .B1(n2100), .C0(n604), 
        .C1(n2103), .Y(n2436) );
  OAI222XL U1741 ( .A0(n652), .A1(n2104), .B0(n644), .B1(n2106), .C0(n636), 
        .C1(n2109), .Y(n2435) );
  OAI222XL U1742 ( .A0(n683), .A1(n2110), .B0(n660), .B1(n2112), .C0(n668), 
        .C1(n2114), .Y(n2434) );
  OAI222XL U1743 ( .A0(n417), .A1(n2117), .B0(n425), .B1(n2118), .C0(n410), 
        .C1(n2120), .Y(n2433) );
  NOR3X1 U1744 ( .A(n2437), .B(n2438), .C(n2439), .Y(n2431) );
  OAI22XL U1745 ( .A0(n516), .A1(n2123), .B0(n500), .B1(n2124), .Y(n2439) );
  OAI22XL U1746 ( .A0(n508), .A1(n2127), .B0(n492), .B1(n2128), .Y(n2438) );
  OAI222XL U1747 ( .A0(n524), .A1(n2130), .B0(n540), .B1(n2132), .C0(n548), 
        .C1(n2135), .Y(n2437) );
  AOI222XL U1748 ( .A0(n2136), .A1(n1706), .B0(n2138), .B1(n1746), .C0(n2384), 
        .C1(n1693), .Y(n2430) );
  AOI222XL U1749 ( .A0(n2143), .A1(n2440), .B0(n2144), .B1(n1722), .C0(n2146), 
        .C1(n1826), .Y(n2429) );
  NAND4X1 U1750 ( .A(n2442), .B(n2443), .C(n2444), .D(n2445), .Y(n2441) );
  NOR4X1 U1751 ( .A(n2446), .B(n2447), .C(n2448), .D(n2449), .Y(n2445) );
  OAI222XL U1752 ( .A0(n619), .A1(n2098), .B0(n611), .B1(n2100), .C0(n603), 
        .C1(n1699), .Y(n2449) );
  OAI222XL U1753 ( .A0(n651), .A1(n2104), .B0(n643), .B1(n2106), .C0(n635), 
        .C1(n2109), .Y(n2448) );
  OAI222XL U1754 ( .A0(n682), .A1(n2110), .B0(n659), .B1(n2112), .C0(n667), 
        .C1(n2114), .Y(n2447) );
  OAI222XL U1755 ( .A0(n416), .A1(n1701), .B0(n424), .B1(n2118), .C0(n409), 
        .C1(n2120), .Y(n2446) );
  NOR3X1 U1756 ( .A(n2450), .B(n2451), .C(n2452), .Y(n2444) );
  OAI22XL U1757 ( .A0(n515), .A1(n1735), .B0(n499), .B1(n2125), .Y(n2452) );
  OAI22XL U1758 ( .A0(n507), .A1(n1736), .B0(n491), .B1(n2128), .Y(n2451) );
  OAI222XL U1759 ( .A0(n523), .A1(n2131), .B0(n539), .B1(n2132), .C0(n547), 
        .C1(n1738), .Y(n2450) );
  AOI222XL U1760 ( .A0(n2136), .A1(n1707), .B0(n2138), .B1(n1747), .C0(n2140), 
        .C1(n1694), .Y(n2443) );
  AOI222XL U1761 ( .A0(n2143), .A1(n2453), .B0(n2144), .B1(n1723), .C0(n2146), 
        .C1(n1827), .Y(n2442) );
  NAND4X1 U1762 ( .A(n2455), .B(n2456), .C(n2457), .D(n2458), .Y(n2454) );
  NOR4X1 U1763 ( .A(n2459), .B(n2460), .C(n2461), .D(n2462), .Y(n2458) );
  OAI222XL U1764 ( .A0(n618), .A1(n2098), .B0(n610), .B1(n2100), .C0(n602), 
        .C1(n2103), .Y(n2462) );
  OAI222XL U1765 ( .A0(n650), .A1(n2104), .B0(n642), .B1(n2106), .C0(n634), 
        .C1(n2109), .Y(n2461) );
  OAI222XL U1766 ( .A0(n681), .A1(n2110), .B0(n658), .B1(n2112), .C0(n666), 
        .C1(n2114), .Y(n2460) );
  OAI222XL U1767 ( .A0(n415), .A1(n2117), .B0(n423), .B1(n2118), .C0(n408), 
        .C1(n2120), .Y(n2459) );
  NOR3X1 U1768 ( .A(n2463), .B(n2464), .C(n2465), .Y(n2457) );
  OAI22XL U1769 ( .A0(n514), .A1(n1735), .B0(n498), .B1(n2124), .Y(n2465) );
  OAI22XL U1770 ( .A0(n506), .A1(n1736), .B0(n490), .B1(n2128), .Y(n2464) );
  OAI222XL U1771 ( .A0(n522), .A1(n2131), .B0(n538), .B1(n2132), .C0(n546), 
        .C1(n1738), .Y(n2463) );
  AOI222XL U1772 ( .A0(n2136), .A1(n1708), .B0(n2138), .B1(n1748), .C0(n2140), 
        .C1(n1695), .Y(n2456) );
  AOI222XL U1773 ( .A0(n2143), .A1(n2466), .B0(n2144), .B1(n1724), .C0(n2146), 
        .C1(n1828), .Y(n2455) );
  NAND4X1 U1774 ( .A(n2468), .B(n2469), .C(n2470), .D(n2471), .Y(n2467) );
  NOR4X1 U1775 ( .A(n2472), .B(n2473), .C(n2474), .D(n2475), .Y(n2471) );
  OAI222XL U1776 ( .A0(n617), .A1(n1741), .B0(n609), .B1(n2100), .C0(n2361), 
        .C1(n2102), .Y(n2475) );
  OAI222XL U1777 ( .A0(n649), .A1(n2104), .B0(n641), .B1(n2106), .C0(n633), 
        .C1(n2109), .Y(n2474) );
  OAI222XL U1778 ( .A0(n2314), .A1(n2110), .B0(n657), .B1(n2112), .C0(n2363), 
        .C1(n2114), .Y(n2473) );
  OAI222XL U1779 ( .A0(n2315), .A1(n2117), .B0(n422), .B1(n2118), .C0(n407), 
        .C1(n2120), .Y(n2472) );
  NOR3X1 U1780 ( .A(n2476), .B(n2477), .C(n2478), .Y(n2470) );
  OAI22XL U1781 ( .A0(n513), .A1(n1735), .B0(n497), .B1(n2380), .Y(n2478) );
  OAI22XL U1782 ( .A0(n505), .A1(n2127), .B0(n489), .B1(n2128), .Y(n2477) );
  OAI222XL U1783 ( .A0(n521), .A1(n2131), .B0(n537), .B1(n2132), .C0(n545), 
        .C1(n1738), .Y(n2476) );
  AOI222XL U1784 ( .A0(n2136), .A1(n1709), .B0(n2138), .B1(n1749), .C0(n2140), 
        .C1(n1696), .Y(n2469) );
  AOI222XL U1785 ( .A0(n2142), .A1(n1773), .B0(n2144), .B1(n1725), .C0(n2146), 
        .C1(n1829), .Y(n2468) );
  NAND4X1 U1786 ( .A(n2480), .B(n2481), .C(n2482), .D(n2483), .Y(n2479) );
  NOR4X1 U1787 ( .A(n2484), .B(n2485), .C(n2486), .D(n2487), .Y(n2483) );
  OAI222XL U1788 ( .A0(n584), .A1(n2099), .B0(n576), .B1(n2100), .C0(n568), 
        .C1(n2103), .Y(n2487) );
  OAI222XL U1789 ( .A0(n616), .A1(n2104), .B0(n608), .B1(n2106), .C0(n600), 
        .C1(n2109), .Y(n2486) );
  OAI222XL U1790 ( .A0(n648), .A1(n2110), .B0(n624), .B1(n2112), .C0(n632), 
        .C1(n2114), .Y(n2485) );
  OAI222XL U1791 ( .A0(n680), .A1(n2117), .B0(n656), .B1(n2118), .C0(n672), 
        .C1(n2120), .Y(n2484) );
  NOR3X1 U1792 ( .A(n2488), .B(n2489), .C(n2490), .Y(n2482) );
  OAI22XL U1793 ( .A0(n480), .A1(n1735), .B0(n464), .B1(n2125), .Y(n2490) );
  OAI22XL U1794 ( .A0(n472), .A1(n2126), .B0(n456), .B1(n2128), .Y(n2489) );
  OAI222XL U1795 ( .A0(n488), .A1(n2131), .B0(n504), .B1(n2132), .C0(n512), 
        .C1(n1738), .Y(n2488) );
  AOI222XL U1796 ( .A0(n2136), .A1(n1806), .B0(n2138), .B1(n1710), .C0(n2140), 
        .C1(n1750), .Y(n2481) );
  AOI222XL U1797 ( .A0(n2143), .A1(n1782), .B0(n2144), .B1(n1689), .C0(n2146), 
        .C1(n1726), .Y(n2480) );
  NAND4X1 U1798 ( .A(n2492), .B(n2493), .C(n2494), .D(n2495), .Y(n2491) );
  NOR4X1 U1799 ( .A(n2496), .B(n2497), .C(n2498), .D(n2499), .Y(n2495) );
  OAI222XL U1800 ( .A0(n583), .A1(n2098), .B0(n575), .B1(n2100), .C0(n567), 
        .C1(n2103), .Y(n2499) );
  OAI222XL U1801 ( .A0(n615), .A1(n2104), .B0(n607), .B1(n2106), .C0(n599), 
        .C1(n2109), .Y(n2498) );
  OAI222XL U1802 ( .A0(n647), .A1(n2110), .B0(n623), .B1(n2112), .C0(n631), 
        .C1(n2114), .Y(n2497) );
  OAI222XL U1803 ( .A0(n679), .A1(n2117), .B0(n655), .B1(n2118), .C0(n671), 
        .C1(n2120), .Y(n2496) );
  NOR3X1 U1804 ( .A(n2500), .B(n2501), .C(n2502), .Y(n2494) );
  OAI22XL U1805 ( .A0(n479), .A1(n1735), .B0(n463), .B1(n2125), .Y(n2502) );
  OAI22XL U1806 ( .A0(n471), .A1(n2127), .B0(n455), .B1(n2128), .Y(n2501) );
  OAI222XL U1807 ( .A0(n487), .A1(n2131), .B0(n503), .B1(n2132), .C0(n511), 
        .C1(n1738), .Y(n2500) );
  AOI222XL U1808 ( .A0(n2136), .A1(n1807), .B0(n2138), .B1(n1711), .C0(n2140), 
        .C1(n1751), .Y(n2493) );
  AOI222XL U1809 ( .A0(n2143), .A1(n1783), .B0(n2144), .B1(n1690), .C0(n2146), 
        .C1(n1727), .Y(n2492) );
  NAND4X1 U1810 ( .A(n2504), .B(n2505), .C(n2506), .D(n2507), .Y(n2503) );
  NOR4X1 U1811 ( .A(n2508), .B(n2509), .C(n2510), .D(n2511), .Y(n2507) );
  OAI222XL U1812 ( .A0(n582), .A1(n2098), .B0(n574), .B1(n2100), .C0(n566), 
        .C1(n2103), .Y(n2511) );
  OAI222XL U1813 ( .A0(n614), .A1(n2104), .B0(n606), .B1(n2106), .C0(n598), 
        .C1(n2109), .Y(n2510) );
  OAI222XL U1814 ( .A0(n646), .A1(n2110), .B0(n622), .B1(n2112), .C0(n630), 
        .C1(n2114), .Y(n2509) );
  OAI222XL U1815 ( .A0(n678), .A1(n2117), .B0(n654), .B1(n2118), .C0(n670), 
        .C1(n2120), .Y(n2508) );
  NOR3X1 U1816 ( .A(n2512), .B(n2513), .C(n2514), .Y(n2506) );
  OAI22XL U1817 ( .A0(n478), .A1(n1735), .B0(n462), .B1(n2125), .Y(n2514) );
  OAI22XL U1818 ( .A0(n470), .A1(n2127), .B0(n454), .B1(n2128), .Y(n2513) );
  OAI222XL U1819 ( .A0(n486), .A1(n2131), .B0(n502), .B1(n2132), .C0(n510), 
        .C1(n1738), .Y(n2512) );
  AOI222XL U1820 ( .A0(n2136), .A1(n1808), .B0(n2138), .B1(n1712), .C0(n2140), 
        .C1(n1752), .Y(n2505) );
  AOI222XL U1821 ( .A0(n2143), .A1(n1784), .B0(n2144), .B1(n1691), .C0(n2146), 
        .C1(n1728), .Y(n2504) );
  NAND4X1 U1822 ( .A(n2516), .B(n2517), .C(n2518), .D(n2519), .Y(n2515) );
  NOR4X1 U1823 ( .A(n2520), .B(n2521), .C(n2522), .D(n2523), .Y(n2519) );
  OAI222XL U1824 ( .A0(n581), .A1(n2098), .B0(n573), .B1(n2100), .C0(n565), 
        .C1(n2103), .Y(n2523) );
  OAI222XL U1825 ( .A0(n613), .A1(n2104), .B0(n605), .B1(n2106), .C0(n597), 
        .C1(n2109), .Y(n2522) );
  OAI222XL U1826 ( .A0(n645), .A1(n2110), .B0(n621), .B1(n2112), .C0(n629), 
        .C1(n2114), .Y(n2521) );
  OAI222XL U1827 ( .A0(n677), .A1(n2117), .B0(n653), .B1(n2118), .C0(n669), 
        .C1(n2120), .Y(n2520) );
  NOR3X1 U1828 ( .A(n2524), .B(n2525), .C(n2526), .Y(n2518) );
  OAI22XL U1829 ( .A0(n477), .A1(n2123), .B0(n461), .B1(n2125), .Y(n2526) );
  OAI22XL U1830 ( .A0(n469), .A1(n2127), .B0(n453), .B1(n2128), .Y(n2525) );
  OAI222XL U1831 ( .A0(n485), .A1(n2131), .B0(n501), .B1(n2132), .C0(n509), 
        .C1(n2135), .Y(n2524) );
  AOI222XL U1832 ( .A0(n2136), .A1(n1809), .B0(n2138), .B1(n1713), .C0(n2140), 
        .C1(n1753), .Y(n2517) );
  AOI222XL U1833 ( .A0(n2143), .A1(n1785), .B0(n2144), .B1(n1692), .C0(n2146), 
        .C1(n1729), .Y(n2516) );
  NAND4X1 U1834 ( .A(n2528), .B(n2529), .C(n2530), .D(n2531), .Y(n2527) );
  NOR4X1 U1835 ( .A(n2532), .B(n2533), .C(n2534), .D(n2535), .Y(n2531) );
  OAI222XL U1836 ( .A0(n580), .A1(n2098), .B0(n572), .B1(n2100), .C0(n564), 
        .C1(n2103), .Y(n2535) );
  OAI222XL U1837 ( .A0(n612), .A1(n2104), .B0(n604), .B1(n2106), .C0(n596), 
        .C1(n2109), .Y(n2534) );
  OAI222XL U1838 ( .A0(n644), .A1(n2111), .B0(n620), .B1(n2112), .C0(n628), 
        .C1(n2114), .Y(n2533) );
  OAI222XL U1839 ( .A0(n676), .A1(n2116), .B0(n652), .B1(n2118), .C0(n668), 
        .C1(n2121), .Y(n2532) );
  NOR3X1 U1840 ( .A(n2536), .B(n2537), .C(n2538), .Y(n2530) );
  OAI22XL U1841 ( .A0(n476), .A1(n2123), .B0(n460), .B1(n2380), .Y(n2538) );
  OAI22XL U1842 ( .A0(n468), .A1(n2127), .B0(n452), .B1(n2128), .Y(n2537) );
  OAI222XL U1843 ( .A0(n484), .A1(n2131), .B0(n500), .B1(n2132), .C0(n508), 
        .C1(n2135), .Y(n2536) );
  AOI222XL U1844 ( .A0(n2137), .A1(n1810), .B0(n2138), .B1(n1714), .C0(n2140), 
        .C1(n1754), .Y(n2529) );
  AOI222XL U1845 ( .A0(n2143), .A1(n1786), .B0(n2145), .B1(n1693), .C0(n2147), 
        .C1(n1730), .Y(n2528) );
  NAND4X1 U1846 ( .A(n2540), .B(n2541), .C(n2542), .D(n2543), .Y(n2539) );
  NOR4X1 U1847 ( .A(n2544), .B(n2545), .C(n2546), .D(n2547), .Y(n2543) );
  OAI222XL U1848 ( .A0(n579), .A1(n2098), .B0(n571), .B1(n2100), .C0(n563), 
        .C1(n1699), .Y(n2547) );
  OAI222XL U1849 ( .A0(n611), .A1(n2105), .B0(n603), .B1(n2107), .C0(n595), 
        .C1(n2109), .Y(n2546) );
  OAI222XL U1850 ( .A0(n643), .A1(n1739), .B0(n619), .B1(n2113), .C0(n627), 
        .C1(n2115), .Y(n2545) );
  OAI222XL U1851 ( .A0(n675), .A1(n2116), .B0(n651), .B1(n2119), .C0(n667), 
        .C1(n1684), .Y(n2544) );
  NOR3X1 U1852 ( .A(n2548), .B(n2549), .C(n2550), .Y(n2542) );
  OAI22XL U1853 ( .A0(n475), .A1(n2123), .B0(n459), .B1(n2125), .Y(n2550) );
  OAI22XL U1854 ( .A0(n467), .A1(n2127), .B0(n451), .B1(n2381), .Y(n2549) );
  OAI222XL U1855 ( .A0(n483), .A1(n2131), .B0(n499), .B1(n2132), .C0(n507), 
        .C1(n2135), .Y(n2548) );
  AOI222XL U1856 ( .A0(n2137), .A1(n1811), .B0(n2139), .B1(n1715), .C0(n2140), 
        .C1(n1755), .Y(n2541) );
  AOI222XL U1857 ( .A0(n2143), .A1(n1787), .B0(n2145), .B1(n1694), .C0(n2147), 
        .C1(n1731), .Y(n2540) );
  NAND4X1 U1858 ( .A(n2552), .B(n2553), .C(n2554), .D(n2555), .Y(n2551) );
  NOR4X1 U1859 ( .A(n2556), .B(n2557), .C(n2558), .D(n2559), .Y(n2555) );
  OAI222XL U1860 ( .A0(n578), .A1(n2098), .B0(n570), .B1(n2100), .C0(n562), 
        .C1(n2103), .Y(n2559) );
  OAI222XL U1861 ( .A0(n610), .A1(n2105), .B0(n602), .B1(n2107), .C0(n594), 
        .C1(n2109), .Y(n2558) );
  OAI222XL U1862 ( .A0(n642), .A1(n2111), .B0(n618), .B1(n2113), .C0(n626), 
        .C1(n2115), .Y(n2557) );
  OAI222XL U1863 ( .A0(n674), .A1(n2116), .B0(n650), .B1(n2119), .C0(n666), 
        .C1(n2121), .Y(n2556) );
  NOR3X1 U1864 ( .A(n2560), .B(n2561), .C(n2562), .Y(n2554) );
  OAI22XL U1865 ( .A0(n474), .A1(n2123), .B0(n458), .B1(n2380), .Y(n2562) );
  OAI22XL U1866 ( .A0(n466), .A1(n2127), .B0(n450), .B1(n2129), .Y(n2561) );
  OAI222XL U1867 ( .A0(n482), .A1(n2131), .B0(n498), .B1(n2132), .C0(n506), 
        .C1(n2135), .Y(n2560) );
  AOI222XL U1868 ( .A0(n2137), .A1(n1812), .B0(n2383), .B1(n1716), .C0(n2140), 
        .C1(n1756), .Y(n2553) );
  AOI222XL U1869 ( .A0(n2143), .A1(n1788), .B0(n2145), .B1(n1695), .C0(n2147), 
        .C1(n1732), .Y(n2552) );
  NAND4X1 U1870 ( .A(n2564), .B(n2565), .C(n2566), .D(n2567), .Y(n2563) );
  NOR4X1 U1871 ( .A(n2568), .B(n2569), .C(n2570), .D(n2571), .Y(n2567) );
  OAI222XL U1872 ( .A0(n577), .A1(n2098), .B0(n569), .B1(n2100), .C0(n561), 
        .C1(n2103), .Y(n2571) );
  OAI222XL U1873 ( .A0(n609), .A1(n2105), .B0(n2361), .B1(n2107), .C0(n593), 
        .C1(n2109), .Y(n2570) );
  OAI222XL U1874 ( .A0(n641), .A1(n2111), .B0(n617), .B1(n2113), .C0(n625), 
        .C1(n2115), .Y(n2569) );
  OAI222XL U1875 ( .A0(n673), .A1(n2116), .B0(n649), .B1(n2119), .C0(n2363), 
        .C1(n2121), .Y(n2568) );
  NOR3X1 U1876 ( .A(n2572), .B(n2573), .C(n2574), .Y(n2566) );
  OAI22XL U1877 ( .A0(n473), .A1(n2123), .B0(n457), .B1(n2125), .Y(n2574) );
  OAI22XL U1878 ( .A0(n465), .A1(n2127), .B0(n449), .B1(n2129), .Y(n2573) );
  OAI222XL U1879 ( .A0(n481), .A1(n2131), .B0(n497), .B1(n2132), .C0(n505), 
        .C1(n2135), .Y(n2572) );
  AOI222XL U1880 ( .A0(n2137), .A1(n1813), .B0(n2138), .B1(n1717), .C0(n2140), 
        .C1(n1757), .Y(n2565) );
  AOI222XL U1881 ( .A0(n2143), .A1(n1789), .B0(n2145), .B1(n1696), .C0(n2147), 
        .C1(n1733), .Y(n2564) );
  NAND4X1 U1882 ( .A(n2576), .B(n2577), .C(n2578), .D(n2579), .Y(n2575) );
  NOR4X1 U1883 ( .A(n2580), .B(n2581), .C(n2582), .D(n2583), .Y(n2579) );
  OAI222XL U1884 ( .A0(n632), .A1(n2098), .B0(n624), .B1(n2100), .C0(n616), 
        .C1(n1699), .Y(n2583) );
  OAI222XL U1885 ( .A0(n664), .A1(n2105), .B0(n656), .B1(n2107), .C0(n648), 
        .C1(n1698), .Y(n2582) );
  OAI222XL U1886 ( .A0(n429), .A1(n1739), .B0(n672), .B1(n2113), .C0(n680), 
        .C1(n2115), .Y(n2581) );
  OAI222XL U1887 ( .A0(n436), .A1(n2116), .B0(n406), .B1(n2119), .C0(n421), 
        .C1(n1684), .Y(n2580) );
  NOR3X1 U1888 ( .A(n2584), .B(n2585), .C(n2586), .Y(n2578) );
  OAI22XL U1889 ( .A0(n528), .A1(n2123), .B0(n512), .B1(n2125), .Y(n2586) );
  OAI22XL U1890 ( .A0(n520), .A1(n2127), .B0(n504), .B1(n2129), .Y(n2585) );
  OAI222XL U1891 ( .A0(n536), .A1(n2131), .B0(n552), .B1(n2132), .C0(n560), 
        .C1(n2135), .Y(n2584) );
  AOI222XL U1892 ( .A0(n2137), .A1(n1814), .B0(n2138), .B1(n1702), .C0(n2140), 
        .C1(n1742), .Y(n2577) );
  AOI222XL U1893 ( .A0(n2143), .A1(n1798), .B0(n2145), .B1(n1766), .C0(n2147), 
        .C1(n1718), .Y(n2576) );
  NAND4X1 U1894 ( .A(n2588), .B(n2589), .C(n2590), .D(n2591), .Y(n2587) );
  NOR4X1 U1895 ( .A(n2592), .B(n2593), .C(n2594), .D(n2595), .Y(n2591) );
  OAI222XL U1896 ( .A0(n631), .A1(n2098), .B0(n623), .B1(n2100), .C0(n615), 
        .C1(n1699), .Y(n2595) );
  OAI222XL U1897 ( .A0(n663), .A1(n2105), .B0(n655), .B1(n2107), .C0(n647), 
        .C1(n1698), .Y(n2594) );
  OAI222XL U1898 ( .A0(n428), .A1(n1739), .B0(n671), .B1(n2113), .C0(n679), 
        .C1(n2115), .Y(n2593) );
  OAI222XL U1899 ( .A0(n435), .A1(n2116), .B0(n405), .B1(n2119), .C0(n420), 
        .C1(n1684), .Y(n2592) );
  NOR3X1 U1900 ( .A(n2596), .B(n2597), .C(n2598), .Y(n2590) );
  OAI22XL U1901 ( .A0(n527), .A1(n2123), .B0(n511), .B1(n2125), .Y(n2598) );
  OAI22XL U1902 ( .A0(n519), .A1(n2127), .B0(n503), .B1(n2129), .Y(n2597) );
  OAI222XL U1903 ( .A0(n535), .A1(n2131), .B0(n551), .B1(n2132), .C0(n559), 
        .C1(n2135), .Y(n2596) );
  AOI222XL U1904 ( .A0(n2137), .A1(n1815), .B0(n2138), .B1(n1703), .C0(n2140), 
        .C1(n1743), .Y(n2589) );
  AOI222XL U1905 ( .A0(n2143), .A1(n1799), .B0(n2145), .B1(n1767), .C0(n2147), 
        .C1(n1719), .Y(n2588) );
  NAND4X1 U1906 ( .A(n2600), .B(n2601), .C(n2602), .D(n2603), .Y(n2599) );
  NOR4X1 U1907 ( .A(n2604), .B(n2605), .C(n2606), .D(n2607), .Y(n2603) );
  OAI222XL U1908 ( .A0(n630), .A1(n2098), .B0(n622), .B1(n2100), .C0(n614), 
        .C1(n2103), .Y(n2607) );
  OAI222XL U1909 ( .A0(n662), .A1(n2105), .B0(n654), .B1(n2107), .C0(n646), 
        .C1(n1698), .Y(n2606) );
  OAI222XL U1910 ( .A0(n427), .A1(n1739), .B0(n670), .B1(n2113), .C0(n678), 
        .C1(n2115), .Y(n2605) );
  OAI222XL U1911 ( .A0(n434), .A1(n2116), .B0(n404), .B1(n2119), .C0(n419), 
        .C1(n2121), .Y(n2604) );
  NOR3X1 U1912 ( .A(n2608), .B(n2609), .C(n2610), .Y(n2602) );
  OAI22XL U1913 ( .A0(n526), .A1(n2123), .B0(n510), .B1(n2380), .Y(n2610) );
  OAI22XL U1914 ( .A0(n518), .A1(n2127), .B0(n502), .B1(n2381), .Y(n2609) );
  OAI222XL U1915 ( .A0(n534), .A1(n2131), .B0(n550), .B1(n2132), .C0(n558), 
        .C1(n2135), .Y(n2608) );
  AOI222XL U1916 ( .A0(n2137), .A1(n1816), .B0(n2383), .B1(n1704), .C0(n2140), 
        .C1(n1744), .Y(n2601) );
  AOI222XL U1917 ( .A0(n2143), .A1(n1800), .B0(n2145), .B1(n1768), .C0(n2147), 
        .C1(n1720), .Y(n2600) );
  NAND4X1 U1918 ( .A(n2612), .B(n2613), .C(n2614), .D(n2615), .Y(n2611) );
  NOR4X1 U1919 ( .A(n2616), .B(n2617), .C(n2618), .D(n2619), .Y(n2615) );
  OAI222XL U1920 ( .A0(n629), .A1(n2098), .B0(n621), .B1(n2100), .C0(n613), 
        .C1(n1699), .Y(n2619) );
  OAI222XL U1921 ( .A0(n661), .A1(n2105), .B0(n653), .B1(n2107), .C0(n645), 
        .C1(n1698), .Y(n2618) );
  OAI222XL U1922 ( .A0(n426), .A1(n1739), .B0(n669), .B1(n2113), .C0(n677), 
        .C1(n2115), .Y(n2617) );
  OAI222XL U1923 ( .A0(n433), .A1(n2116), .B0(n403), .B1(n2119), .C0(n418), 
        .C1(n1684), .Y(n2616) );
  NOR3X1 U1924 ( .A(n2620), .B(n2621), .C(n2622), .Y(n2614) );
  OAI22XL U1925 ( .A0(n525), .A1(n2123), .B0(n509), .B1(n2125), .Y(n2622) );
  OAI22XL U1926 ( .A0(n517), .A1(n2127), .B0(n501), .B1(n2381), .Y(n2621) );
  OAI222XL U1927 ( .A0(n533), .A1(n2131), .B0(n549), .B1(n2132), .C0(n557), 
        .C1(n2135), .Y(n2620) );
  AOI222XL U1928 ( .A0(n2137), .A1(n1817), .B0(n2138), .B1(n1705), .C0(n2140), 
        .C1(n1745), .Y(n2613) );
  AOI222XL U1929 ( .A0(n2143), .A1(n1801), .B0(n2145), .B1(n1769), .C0(n2147), 
        .C1(n1721), .Y(n2612) );
  NAND4X1 U1930 ( .A(n2624), .B(n2625), .C(n2626), .D(n2627), .Y(n2623) );
  NOR4X1 U1931 ( .A(n2628), .B(n2629), .C(n2630), .D(n2631), .Y(n2627) );
  OAI222XL U1932 ( .A0(n628), .A1(n2098), .B0(n620), .B1(n2100), .C0(n612), 
        .C1(n2103), .Y(n2631) );
  OAI222XL U1933 ( .A0(n660), .A1(n2105), .B0(n652), .B1(n2107), .C0(n644), 
        .C1(n2109), .Y(n2630) );
  OAI222XL U1934 ( .A0(n425), .A1(n2111), .B0(n668), .B1(n2113), .C0(n676), 
        .C1(n2115), .Y(n2629) );
  OAI222XL U1935 ( .A0(n432), .A1(n2116), .B0(n402), .B1(n2119), .C0(n417), 
        .C1(n2121), .Y(n2628) );
  NOR3X1 U1936 ( .A(n2632), .B(n2633), .C(n2634), .Y(n2626) );
  OAI22XL U1937 ( .A0(n524), .A1(n2123), .B0(n508), .B1(n2125), .Y(n2634) );
  OAI22XL U1938 ( .A0(n516), .A1(n2127), .B0(n500), .B1(n2381), .Y(n2633) );
  OAI222XL U1939 ( .A0(n532), .A1(n2131), .B0(n548), .B1(n2132), .C0(n556), 
        .C1(n2135), .Y(n2632) );
  AOI222XL U1940 ( .A0(n2137), .A1(n1818), .B0(n2383), .B1(n1706), .C0(n2140), 
        .C1(n1746), .Y(n2625) );
  AOI222XL U1941 ( .A0(n2142), .A1(n1802), .B0(n2145), .B1(n1770), .C0(n2147), 
        .C1(n1722), .Y(n2624) );
  NAND4X1 U1942 ( .A(n2636), .B(n2637), .C(n2638), .D(n2639), .Y(n2635) );
  NOR4X1 U1943 ( .A(n2640), .B(n2641), .C(n2642), .D(n2643), .Y(n2639) );
  OAI222XL U1944 ( .A0(n627), .A1(n2098), .B0(n619), .B1(n2100), .C0(n611), 
        .C1(n2103), .Y(n2643) );
  OAI222XL U1945 ( .A0(n659), .A1(n2105), .B0(n651), .B1(n2107), .C0(n643), 
        .C1(n1698), .Y(n2642) );
  OAI222XL U1946 ( .A0(n424), .A1(n2111), .B0(n667), .B1(n2113), .C0(n675), 
        .C1(n2115), .Y(n2641) );
  OAI222XL U1947 ( .A0(n431), .A1(n2116), .B0(n401), .B1(n2119), .C0(n416), 
        .C1(n1684), .Y(n2640) );
  NOR3X1 U1948 ( .A(n2644), .B(n2645), .C(n2646), .Y(n2638) );
  OAI22XL U1949 ( .A0(n523), .A1(n2123), .B0(n507), .B1(n2125), .Y(n2646) );
  OAI22XL U1950 ( .A0(n515), .A1(n2127), .B0(n499), .B1(n2381), .Y(n2645) );
  OAI222XL U1951 ( .A0(n531), .A1(n2131), .B0(n547), .B1(n2132), .C0(n555), 
        .C1(n2135), .Y(n2644) );
  AOI222XL U1952 ( .A0(n2137), .A1(n1819), .B0(n2138), .B1(n1707), .C0(n2140), 
        .C1(n1747), .Y(n2637) );
  AOI222XL U1953 ( .A0(n2142), .A1(n1803), .B0(n2145), .B1(n1771), .C0(n2147), 
        .C1(n1723), .Y(n2636) );
  NAND4X1 U1954 ( .A(n2648), .B(n2649), .C(n2650), .D(n2651), .Y(n2647) );
  NOR4X1 U1955 ( .A(n2652), .B(n2653), .C(n2654), .D(n2655), .Y(n2651) );
  OAI222XL U1956 ( .A0(n626), .A1(n2098), .B0(n618), .B1(n2100), .C0(n610), 
        .C1(n2103), .Y(n2655) );
  OAI222XL U1957 ( .A0(n658), .A1(n2105), .B0(n650), .B1(n2107), .C0(n642), 
        .C1(n1698), .Y(n2654) );
  OAI222XL U1958 ( .A0(n423), .A1(n2111), .B0(n666), .B1(n2113), .C0(n674), 
        .C1(n2115), .Y(n2653) );
  OAI222XL U1959 ( .A0(n430), .A1(n2116), .B0(n400), .B1(n2119), .C0(n415), 
        .C1(n1684), .Y(n2652) );
  NOR3X1 U1960 ( .A(n2656), .B(n2657), .C(n2658), .Y(n2650) );
  OAI22XL U1961 ( .A0(n522), .A1(n2123), .B0(n506), .B1(n2125), .Y(n2658) );
  OAI22XL U1962 ( .A0(n514), .A1(n2127), .B0(n498), .B1(n2381), .Y(n2657) );
  OAI222XL U1963 ( .A0(n530), .A1(n2131), .B0(n546), .B1(n2132), .C0(n554), 
        .C1(n2135), .Y(n2656) );
  AOI222XL U1964 ( .A0(n2137), .A1(n1820), .B0(n2138), .B1(n1708), .C0(n2140), 
        .C1(n1748), .Y(n2649) );
  AOI222XL U1965 ( .A0(n2142), .A1(n1804), .B0(n2145), .B1(n1772), .C0(n2147), 
        .C1(n1724), .Y(n2648) );
  NAND4X1 U1966 ( .A(n2660), .B(n2661), .C(n2662), .D(n2663), .Y(n2659) );
  NOR4X1 U1967 ( .A(n2664), .B(n2665), .C(n2666), .D(n2667), .Y(n2663) );
  OAI222XL U1968 ( .A0(n625), .A1(n2099), .B0(n617), .B1(n2101), .C0(n609), 
        .C1(n2102), .Y(n2667) );
  OAI222XL U1969 ( .A0(n657), .A1(n2105), .B0(n649), .B1(n2107), .C0(n641), 
        .C1(n2108), .Y(n2666) );
  OAI222XL U1970 ( .A0(n422), .A1(n1739), .B0(n2363), .B1(n2113), .C0(n673), 
        .C1(n2115), .Y(n2665) );
  OAI222XL U1971 ( .A0(n2313), .A1(n2116), .B0(n399), .B1(n2119), .C0(n2315), 
        .C1(n2121), .Y(n2664) );
  NOR3X1 U1972 ( .A(n2668), .B(n2669), .C(n2670), .Y(n2662) );
  OAI22XL U1973 ( .A0(n521), .A1(n2122), .B0(n505), .B1(n2125), .Y(n2670) );
  OAI22XL U1974 ( .A0(n513), .A1(n2126), .B0(n497), .B1(n2129), .Y(n2669) );
  OAI222XL U1975 ( .A0(n529), .A1(n2130), .B0(n545), .B1(n2133), .C0(n553), 
        .C1(n2134), .Y(n2668) );
  AOI222XL U1976 ( .A0(n2137), .A1(n1821), .B0(n2138), .B1(n1709), .C0(n2141), 
        .C1(n1749), .Y(n2661) );
  AOI222XL U1977 ( .A0(n2142), .A1(n1805), .B0(n2145), .B1(m43_7_), .C0(n2147), 
        .C1(n1725), .Y(n2660) );
  NAND3X1 U1978 ( .A(n2118), .B(n1701), .C(n2676), .Y(n2675) );
  NAND3X1 U1979 ( .A(n2112), .B(n2110), .C(n2120), .Y(n2674) );
  NAND4X1 U1980 ( .A(n2106), .B(n2104), .C(n2114), .D(n2677), .Y(n2673) );
  AND4X1 U1981 ( .A(n2102), .B(n2099), .C(n2101), .D(n2108), .Y(n2677) );
  NAND4X1 U1982 ( .A(n2678), .B(n2679), .C(n2680), .D(n2681), .Y(n2672) );
  NOR3X1 U1983 ( .A(n2136), .B(n2146), .C(n2144), .Y(n2681) );
  NOR3BXL U1984 ( .AN(n2134), .B(n2141), .C(n2139), .Y(n2680) );
  AND3X1 U1985 ( .A(n2122), .B(n1700), .C(n2133), .Y(n2679) );
  AND3X1 U1986 ( .A(n2129), .B(n2124), .C(n2126), .Y(n2678) );
  CLKINVX1 U1987 ( .A(n2682), .Y(n2671) );
  AO22X1 U1988 ( .A0(t11[0]), .A1(n2089), .B0(n2684), .B1(n2685), .Y(n1621) );
  NAND4X1 U1989 ( .A(n2686), .B(n2687), .C(n2688), .D(n2689), .Y(n2685) );
  NOR4X1 U1990 ( .A(n2690), .B(n2691), .C(n2692), .D(n2693), .Y(n2689) );
  OAI222XL U1991 ( .A0(n576), .A1(n2099), .B0(n568), .B1(n2101), .C0(n560), 
        .C1(n2102), .Y(n2693) );
  OAI222XL U1992 ( .A0(n608), .A1(n2105), .B0(n600), .B1(n2107), .C0(n592), 
        .C1(n2108), .Y(n2692) );
  OAI222XL U1993 ( .A0(n640), .A1(n2111), .B0(n616), .B1(n2113), .C0(n624), 
        .C1(n2115), .Y(n2691) );
  OAI222XL U1994 ( .A0(n672), .A1(n2116), .B0(n648), .B1(n2119), .C0(n664), 
        .C1(n2121), .Y(n2690) );
  NOR3X1 U1995 ( .A(n2694), .B(n2695), .C(n2696), .Y(n2688) );
  OAI22XL U1996 ( .A0(n472), .A1(n2122), .B0(n456), .B1(n2124), .Y(n2696) );
  OAI22XL U1997 ( .A0(n464), .A1(n2126), .B0(n448), .B1(n2129), .Y(n2695) );
  OAI222XL U1998 ( .A0(n480), .A1(n2130), .B0(n496), .B1(n2133), .C0(n504), 
        .C1(n2134), .Y(n2694) );
  AOI222XL U1999 ( .A0(n2137), .A1(n1710), .B0(n2139), .B1(n1750), .C0(n2141), 
        .C1(n1790), .Y(n2687) );
  AOI222XL U2000 ( .A0(n2142), .A1(n1758), .B0(n2145), .B1(n1726), .C0(n2147), 
        .C1(n1830), .Y(n2686) );
  AO22X1 U2001 ( .A0(t11[1]), .A1(n2089), .B0(n2684), .B1(n2697), .Y(n1620) );
  NAND4X1 U2002 ( .A(n2698), .B(n2699), .C(n2700), .D(n2701), .Y(n2697) );
  NOR4X1 U2003 ( .A(n2702), .B(n2703), .C(n2704), .D(n2705), .Y(n2701) );
  OAI222XL U2004 ( .A0(n575), .A1(n2099), .B0(n567), .B1(n2101), .C0(n559), 
        .C1(n2102), .Y(n2705) );
  OAI222XL U2005 ( .A0(n607), .A1(n2105), .B0(n599), .B1(n2107), .C0(n591), 
        .C1(n2108), .Y(n2704) );
  OAI222XL U2006 ( .A0(n639), .A1(n2111), .B0(n615), .B1(n2113), .C0(n623), 
        .C1(n2115), .Y(n2703) );
  OAI222XL U2007 ( .A0(n671), .A1(n2116), .B0(n647), .B1(n2119), .C0(n663), 
        .C1(n2121), .Y(n2702) );
  NOR3X1 U2008 ( .A(n2706), .B(n2707), .C(n2708), .Y(n2700) );
  OAI22XL U2009 ( .A0(n471), .A1(n2122), .B0(n455), .B1(n2124), .Y(n2708) );
  OAI22XL U2010 ( .A0(n463), .A1(n2126), .B0(n447), .B1(n2129), .Y(n2707) );
  OAI222XL U2011 ( .A0(n479), .A1(n2130), .B0(n495), .B1(n2133), .C0(n503), 
        .C1(n2134), .Y(n2706) );
  AOI222XL U2012 ( .A0(n2137), .A1(n1711), .B0(n2139), .B1(n1751), .C0(n2141), 
        .C1(n1791), .Y(n2699) );
  AOI222XL U2013 ( .A0(n2142), .A1(n1759), .B0(n2145), .B1(n1727), .C0(n2147), 
        .C1(n1831), .Y(n2698) );
  AO22X1 U2014 ( .A0(t11[2]), .A1(n2089), .B0(n2684), .B1(n2709), .Y(n1619) );
  NAND4X1 U2015 ( .A(n2710), .B(n2711), .C(n2712), .D(n2713), .Y(n2709) );
  NOR4X1 U2016 ( .A(n2714), .B(n2715), .C(n2716), .D(n2717), .Y(n2713) );
  OAI222XL U2017 ( .A0(n574), .A1(n2099), .B0(n566), .B1(n2101), .C0(n558), 
        .C1(n2102), .Y(n2717) );
  OAI222XL U2018 ( .A0(n606), .A1(n2105), .B0(n598), .B1(n1737), .C0(n590), 
        .C1(n2108), .Y(n2716) );
  OAI222XL U2019 ( .A0(n638), .A1(n2111), .B0(n614), .B1(n2113), .C0(n622), 
        .C1(n2115), .Y(n2715) );
  OAI222XL U2020 ( .A0(n670), .A1(n2117), .B0(n646), .B1(n2119), .C0(n662), 
        .C1(n2121), .Y(n2714) );
  NOR3X1 U2021 ( .A(n2718), .B(n2719), .C(n2720), .Y(n2712) );
  OAI22XL U2022 ( .A0(n470), .A1(n2122), .B0(n454), .B1(n2124), .Y(n2720) );
  OAI22XL U2023 ( .A0(n462), .A1(n2126), .B0(n446), .B1(n2129), .Y(n2719) );
  OAI222XL U2024 ( .A0(n478), .A1(n2130), .B0(n494), .B1(n2133), .C0(n502), 
        .C1(n2134), .Y(n2718) );
  AOI222XL U2025 ( .A0(n2137), .A1(n1712), .B0(n2139), .B1(n1752), .C0(n2141), 
        .C1(n1792), .Y(n2711) );
  AOI222XL U2026 ( .A0(n2142), .A1(n1760), .B0(n2145), .B1(n1728), .C0(n2147), 
        .C1(n1832), .Y(n2710) );
  AO22X1 U2027 ( .A0(t11[3]), .A1(n2089), .B0(n2684), .B1(n2721), .Y(n1618) );
  NAND4X1 U2028 ( .A(n2722), .B(n2723), .C(n2724), .D(n2725), .Y(n2721) );
  NOR4X1 U2029 ( .A(n2726), .B(n2727), .C(n2728), .D(n2729), .Y(n2725) );
  OAI222XL U2030 ( .A0(n573), .A1(n2099), .B0(n565), .B1(n2101), .C0(n557), 
        .C1(n2102), .Y(n2729) );
  OAI222XL U2031 ( .A0(n605), .A1(n2105), .B0(n597), .B1(n1737), .C0(n589), 
        .C1(n2108), .Y(n2728) );
  OAI222XL U2032 ( .A0(n637), .A1(n2111), .B0(n613), .B1(n2113), .C0(n621), 
        .C1(n2115), .Y(n2727) );
  OAI222XL U2033 ( .A0(n669), .A1(n2117), .B0(n645), .B1(n2119), .C0(n661), 
        .C1(n2121), .Y(n2726) );
  NOR3X1 U2034 ( .A(n2730), .B(n2731), .C(n2732), .Y(n2724) );
  OAI22XL U2035 ( .A0(n469), .A1(n2122), .B0(n453), .B1(n2124), .Y(n2732) );
  OAI22XL U2036 ( .A0(n461), .A1(n2126), .B0(n445), .B1(n2129), .Y(n2731) );
  OAI222XL U2037 ( .A0(n477), .A1(n2130), .B0(n493), .B1(n2133), .C0(n501), 
        .C1(n2134), .Y(n2730) );
  AOI222XL U2038 ( .A0(n2137), .A1(n1713), .B0(n2139), .B1(n1753), .C0(n2141), 
        .C1(n1793), .Y(n2723) );
  AOI222XL U2039 ( .A0(n2142), .A1(n1761), .B0(n2145), .B1(n1729), .C0(n2147), 
        .C1(n1833), .Y(n2722) );
  AO22X1 U2040 ( .A0(t11[4]), .A1(n2089), .B0(n2684), .B1(n2733), .Y(n1617) );
  NAND4X1 U2041 ( .A(n2734), .B(n2735), .C(n2736), .D(n2737), .Y(n2733) );
  NOR4X1 U2042 ( .A(n2738), .B(n2739), .C(n2740), .D(n2741), .Y(n2737) );
  OAI222XL U2043 ( .A0(n572), .A1(n2099), .B0(n564), .B1(n2101), .C0(n556), 
        .C1(n2102), .Y(n2741) );
  OAI222XL U2044 ( .A0(n604), .A1(n2105), .B0(n596), .B1(n1737), .C0(n588), 
        .C1(n2108), .Y(n2740) );
  OAI222XL U2045 ( .A0(n636), .A1(n2111), .B0(n612), .B1(n2113), .C0(n620), 
        .C1(n2115), .Y(n2739) );
  OAI222XL U2046 ( .A0(n668), .A1(n2117), .B0(n644), .B1(n2119), .C0(n660), 
        .C1(n2121), .Y(n2738) );
  NOR3X1 U2047 ( .A(n2742), .B(n2743), .C(n2744), .Y(n2736) );
  OAI22XL U2048 ( .A0(n468), .A1(n2122), .B0(n452), .B1(n2124), .Y(n2744) );
  OAI22XL U2049 ( .A0(n460), .A1(n2126), .B0(n444), .B1(n2129), .Y(n2743) );
  OAI222XL U2050 ( .A0(n476), .A1(n2130), .B0(n492), .B1(n2133), .C0(n500), 
        .C1(n2134), .Y(n2742) );
  AOI222XL U2051 ( .A0(n2137), .A1(n1714), .B0(n2139), .B1(n1754), .C0(n2141), 
        .C1(n1794), .Y(n2735) );
  AOI222XL U2052 ( .A0(n2142), .A1(n1762), .B0(n2145), .B1(n1730), .C0(n2147), 
        .C1(n1834), .Y(n2734) );
  AO22X1 U2053 ( .A0(t11[5]), .A1(n2089), .B0(n2684), .B1(n2745), .Y(n1616) );
  NAND4X1 U2054 ( .A(n2746), .B(n2747), .C(n2748), .D(n2749), .Y(n2745) );
  NOR4X1 U2055 ( .A(n2750), .B(n2751), .C(n2752), .D(n2753), .Y(n2749) );
  OAI222XL U2056 ( .A0(n571), .A1(n2099), .B0(n563), .B1(n2101), .C0(n555), 
        .C1(n2102), .Y(n2753) );
  OAI222XL U2057 ( .A0(n603), .A1(n2105), .B0(n595), .B1(n1737), .C0(n587), 
        .C1(n2108), .Y(n2752) );
  OAI222XL U2058 ( .A0(n635), .A1(n2111), .B0(n611), .B1(n2113), .C0(n619), 
        .C1(n2115), .Y(n2751) );
  OAI222XL U2059 ( .A0(n667), .A1(n2117), .B0(n643), .B1(n2119), .C0(n659), 
        .C1(n2121), .Y(n2750) );
  NOR3X1 U2060 ( .A(n2754), .B(n2755), .C(n2756), .Y(n2748) );
  OAI22XL U2061 ( .A0(n467), .A1(n2122), .B0(n451), .B1(n2124), .Y(n2756) );
  OAI22XL U2062 ( .A0(n459), .A1(n2126), .B0(n443), .B1(n2129), .Y(n2755) );
  OAI222XL U2063 ( .A0(n475), .A1(n2130), .B0(n491), .B1(n2133), .C0(n499), 
        .C1(n2134), .Y(n2754) );
  AOI222XL U2064 ( .A0(n2137), .A1(n1715), .B0(n2139), .B1(n1755), .C0(n2141), 
        .C1(n1795), .Y(n2747) );
  AOI222XL U2065 ( .A0(n2142), .A1(n1763), .B0(n2145), .B1(n1731), .C0(n2147), 
        .C1(n1835), .Y(n2746) );
  AO22X1 U2066 ( .A0(t11[6]), .A1(n2089), .B0(n2684), .B1(n2757), .Y(n1615) );
  NAND4X1 U2067 ( .A(n2758), .B(n2759), .C(n2760), .D(n2761), .Y(n2757) );
  NOR4X1 U2068 ( .A(n2762), .B(n2763), .C(n2764), .D(n2765), .Y(n2761) );
  OAI222XL U2069 ( .A0(n570), .A1(n2099), .B0(n562), .B1(n2101), .C0(n554), 
        .C1(n2102), .Y(n2765) );
  OAI222XL U2070 ( .A0(n602), .A1(n2105), .B0(n594), .B1(n2107), .C0(n586), 
        .C1(n2108), .Y(n2764) );
  OAI222XL U2071 ( .A0(n634), .A1(n2111), .B0(n610), .B1(n2113), .C0(n618), 
        .C1(n2115), .Y(n2763) );
  OAI222XL U2072 ( .A0(n666), .A1(n2117), .B0(n642), .B1(n2119), .C0(n658), 
        .C1(n2121), .Y(n2762) );
  NOR3X1 U2073 ( .A(n2766), .B(n2767), .C(n2768), .Y(n2760) );
  OAI22XL U2074 ( .A0(n466), .A1(n2122), .B0(n450), .B1(n2125), .Y(n2768) );
  OAI22XL U2075 ( .A0(n458), .A1(n2126), .B0(n442), .B1(n2129), .Y(n2767) );
  OAI222XL U2076 ( .A0(n474), .A1(n2130), .B0(n490), .B1(n2133), .C0(n498), 
        .C1(n2134), .Y(n2766) );
  AOI222XL U2077 ( .A0(n2137), .A1(n1716), .B0(n2383), .B1(n1756), .C0(n2141), 
        .C1(n1796), .Y(n2759) );
  AOI222XL U2078 ( .A0(n2142), .A1(n1764), .B0(n2145), .B1(n1732), .C0(n2147), 
        .C1(n1836), .Y(n2758) );
  AO22X1 U2079 ( .A0(t11[7]), .A1(n2089), .B0(n2684), .B1(n2769), .Y(n1614) );
  NAND4X1 U2080 ( .A(n2770), .B(n2771), .C(n2772), .D(n2773), .Y(n2769) );
  NOR4X1 U2081 ( .A(n2774), .B(n2775), .C(n2776), .D(n2777), .Y(n2773) );
  OAI222XL U2082 ( .A0(n569), .A1(n1741), .B0(n561), .B1(n1683), .C0(n553), 
        .C1(n2103), .Y(n2777) );
  OAI222XL U2083 ( .A0(n2361), .A1(n2104), .B0(n593), .B1(n2106), .C0(n585), 
        .C1(n2109), .Y(n2776) );
  CLKINVX1 U2084 ( .A(m43_7_), .Y(n2361) );
  OAI222XL U2085 ( .A0(n633), .A1(n2110), .B0(n609), .B1(n2112), .C0(n617), 
        .C1(n2114), .Y(n2775) );
  OAI222XL U2086 ( .A0(n2363), .A1(n1701), .B0(n641), .B1(n2118), .C0(n657), 
        .C1(n2120), .Y(n2774) );
  CLKINVX1 U2087 ( .A(m55_7_), .Y(n2363) );
  NOR3X1 U2088 ( .A(n2786), .B(n2787), .C(n2788), .Y(n2772) );
  OAI22XL U2089 ( .A0(n465), .A1(n2123), .B0(n449), .B1(n2380), .Y(n2788) );
  OAI22XL U2090 ( .A0(n457), .A1(n2127), .B0(n441), .B1(n2128), .Y(n2787) );
  OAI222XL U2091 ( .A0(n473), .A1(n2130), .B0(n489), .B1(n1685), .C0(n497), 
        .C1(n2135), .Y(n2786) );
  CLKINVX1 U2092 ( .A(n2790), .Y(n2780) );
  CLKINVX1 U2093 ( .A(n2791), .Y(n2779) );
  AND2X1 U2094 ( .A(n2792), .B(n2317), .Y(n2789) );
  AOI222XL U2095 ( .A0(n2136), .A1(n1717), .B0(n2138), .B1(n1757), .C0(n2141), 
        .C1(n1797), .Y(n2771) );
  AND2X1 U2096 ( .A(n2778), .B(n2783), .Y(n2383) );
  AND2X1 U2097 ( .A(n2778), .B(n2354), .Y(n2382) );
  CLKINVX1 U2098 ( .A(n2793), .Y(n2354) );
  AOI222XL U2099 ( .A0(n2142), .A1(n1765), .B0(n2144), .B1(n1733), .C0(n2146), 
        .C1(n1837), .Y(n2770) );
  AND2X1 U2100 ( .A(n2778), .B(n2357), .Y(n2388) );
  CLKINVX1 U2101 ( .A(n2794), .Y(n2357) );
  AND2X1 U2102 ( .A(n2778), .B(n2359), .Y(n2387) );
  CLKINVX1 U2103 ( .A(n2795), .Y(n2359) );
  CLKINVX1 U2104 ( .A(n2676), .Y(n2385) );
  NAND2X1 U2105 ( .A(n2782), .B(n2781), .Y(n2676) );
  CLKINVX1 U2106 ( .A(n2797), .Y(n2781) );
  NOR3X1 U2107 ( .A(n383), .B(n385), .C(n2785), .Y(n2796) );
  OAI31XL U2108 ( .A0(n2799), .A1(start_1_), .A2(n398), .B0(n2172), .Y(n2798)
         );
  AOI31X1 U2109 ( .A0(n2800), .A1(mode[5]), .A2(n2801), .B0(n2802), .Y(n2799)
         );
  NOR4X1 U2110 ( .A(n2317), .B(n2803), .C(mode[7]), .D(n2804), .Y(n2802) );
  OAI21XL U2111 ( .A0(n386), .A1(n2351), .B0(n385), .Y(n2800) );
  AO22X1 U2112 ( .A0(node[0]), .A1(n2805), .B0(N1001), .B1(n2806), .Y(n1613)
         );
  AO22X1 U2113 ( .A0(node[1]), .A1(n2805), .B0(N1002), .B1(n2806), .Y(n1612)
         );
  AO22X1 U2114 ( .A0(node[2]), .A1(n2805), .B0(N1003), .B1(n2806), .Y(n1611)
         );
  AO22X1 U2115 ( .A0(node[3]), .A1(n2805), .B0(N1004), .B1(n2806), .Y(n1610)
         );
  AO22X1 U2116 ( .A0(node[4]), .A1(n2805), .B0(N1005), .B1(n2806), .Y(n1609)
         );
  AO22X1 U2117 ( .A0(node[5]), .A1(n2805), .B0(N1006), .B1(n2806), .Y(n1608)
         );
  AO22X1 U2118 ( .A0(node[6]), .A1(n2805), .B0(N1007), .B1(n2806), .Y(n1607)
         );
  AO22X1 U2119 ( .A0(node[7]), .A1(n2805), .B0(N1008), .B1(n2806), .Y(n1606)
         );
  OAI221XL U2120 ( .A0(n2809), .A1(n2148), .B0(n2149), .B1(n2181), .C0(n2172), 
        .Y(n1604) );
  OAI221XL U2121 ( .A0(n2810), .A1(n2148), .B0(n2149), .B1(n2182), .C0(n2172), 
        .Y(n1603) );
  OAI221XL U2122 ( .A0(n2811), .A1(n2148), .B0(n2149), .B1(n2183), .C0(n2171), 
        .Y(n1602) );
  OAI221XL U2123 ( .A0(n2812), .A1(n2148), .B0(n2149), .B1(n2184), .C0(n2172), 
        .Y(n1601) );
  OAI221XL U2124 ( .A0(n2813), .A1(n2148), .B0(n2149), .B1(n2185), .C0(n2172), 
        .Y(n1600) );
  OAI221XL U2125 ( .A0(n2814), .A1(n2148), .B0(n2149), .B1(n2186), .C0(n2172), 
        .Y(n1599) );
  OAI221XL U2126 ( .A0(n2815), .A1(n2148), .B0(n2149), .B1(n2187), .C0(n2172), 
        .Y(n1598) );
  OAI221XL U2127 ( .A0(n2818), .A1(n2148), .B0(n2149), .B1(n2188), .C0(n2171), 
        .Y(n1596) );
  OAI221XL U2128 ( .A0(n2819), .A1(n2148), .B0(n2149), .B1(n2189), .C0(n2171), 
        .Y(n1595) );
  OAI221XL U2129 ( .A0(n2820), .A1(n2148), .B0(n2149), .B1(n2190), .C0(n2171), 
        .Y(n1594) );
  OAI221XL U2130 ( .A0(n2821), .A1(n2148), .B0(n2149), .B1(n2191), .C0(n2171), 
        .Y(n1593) );
  OAI221XL U2131 ( .A0(n2822), .A1(n2148), .B0(n2149), .B1(n2192), .C0(n2171), 
        .Y(n1592) );
  OAI221XL U2132 ( .A0(n2823), .A1(n2148), .B0(n2149), .B1(n2193), .C0(n2171), 
        .Y(n1591) );
  OAI221XL U2133 ( .A0(n2824), .A1(n2148), .B0(n2149), .B1(n2194), .C0(n2171), 
        .Y(n1590) );
  OAI221XL U2134 ( .A0(n2826), .A1(n2148), .B0(n1949), .B1(n2196), .C0(n2171), 
        .Y(n1588) );
  OAI221XL U2135 ( .A0(n2827), .A1(n2148), .B0(n1949), .B1(n2197), .C0(n2171), 
        .Y(n1587) );
  OAI221XL U2136 ( .A0(n2828), .A1(n2148), .B0(n1949), .B1(n2198), .C0(n2171), 
        .Y(n1586) );
  OAI221XL U2137 ( .A0(n2829), .A1(n2148), .B0(n2149), .B1(n2199), .C0(n2171), 
        .Y(n1585) );
  OAI221XL U2138 ( .A0(n2830), .A1(n2148), .B0(n2149), .B1(n2200), .C0(n2171), 
        .Y(n1584) );
  OAI221XL U2139 ( .A0(n2831), .A1(n2148), .B0(n2149), .B1(n2201), .C0(n2171), 
        .Y(n1583) );
  OAI221XL U2140 ( .A0(n2833), .A1(n2148), .B0(n2149), .B1(n2203), .C0(n2173), 
        .Y(n1581) );
  OAI221XL U2141 ( .A0(n2834), .A1(n2148), .B0(n2149), .B1(n2204), .C0(n2173), 
        .Y(n1580) );
  OAI221XL U2142 ( .A0(n2835), .A1(n2148), .B0(n2149), .B1(n2205), .C0(n2171), 
        .Y(n1579) );
  OAI221XL U2143 ( .A0(n2836), .A1(n2148), .B0(n2149), .B1(n2206), .C0(n2171), 
        .Y(n1578) );
  OAI221XL U2144 ( .A0(n2837), .A1(n2148), .B0(n2149), .B1(n2207), .C0(n2171), 
        .Y(n1577) );
  OAI221XL U2145 ( .A0(n2838), .A1(n2148), .B0(n1949), .B1(n2208), .C0(n2171), 
        .Y(n1576) );
  OAI221XL U2146 ( .A0(n2839), .A1(n2148), .B0(n1949), .B1(n2209), .C0(n2173), 
        .Y(n1575) );
  OAI22XL U2147 ( .A0(n2149), .A1(n2842), .B0(N858), .B1(n2148), .Y(n1572) );
  OAI22XL U2148 ( .A0(n2149), .A1(n2843), .B0(N885), .B1(n2148), .Y(n1571) );
  OAI22XL U2149 ( .A0(n2149), .A1(n2844), .B0(n2088), .B1(n2148), .Y(n1570) );
  OAI21XL U2150 ( .A0(n2847), .A1(n2848), .B0(n2323), .Y(n2846) );
  CLKINVX1 U2151 ( .A(n2849), .Y(n2848) );
  AOI211X1 U2152 ( .A0(n2850), .A1(n2851), .B0(n2852), .C0(n2321), .Y(n2849)
         );
  OAI211X1 U2153 ( .A0(n2853), .A1(n2854), .B0(n2855), .C0(n2856), .Y(n2321)
         );
  NAND2X1 U2154 ( .A(node[3]), .B(n2857), .Y(n2854) );
  NAND3X1 U2155 ( .A(n2858), .B(n2859), .C(n2860), .Y(n2847) );
  CLKINVX1 U2156 ( .A(a2[1]), .Y(n2845) );
  OAI21XL U2157 ( .A0(n2320), .A1(n2861), .B0(n2862), .Y(n1568) );
  CLKINVX1 U2158 ( .A(a2[2]), .Y(n2861) );
  OAI21XL U2159 ( .A0(n2320), .A1(n2863), .B0(n2862), .Y(n1567) );
  CLKINVX1 U2160 ( .A(a2[3]), .Y(n2863) );
  OAI21XL U2161 ( .A0(n2320), .A1(n2864), .B0(n2862), .Y(n1566) );
  CLKINVX1 U2162 ( .A(a2[4]), .Y(n2864) );
  OAI21XL U2163 ( .A0(n2320), .A1(n2865), .B0(n2862), .Y(n1565) );
  CLKINVX1 U2164 ( .A(a2[5]), .Y(n2865) );
  OAI21XL U2165 ( .A0(n2320), .A1(n2866), .B0(n2862), .Y(n1564) );
  CLKINVX1 U2166 ( .A(a2[6]), .Y(n2866) );
  OAI21XL U2167 ( .A0(n2320), .A1(n2867), .B0(n2862), .Y(n1563) );
  CLKINVX1 U2168 ( .A(a2[7]), .Y(n2867) );
  OAI21XL U2169 ( .A0(n2320), .A1(n2868), .B0(n2862), .Y(n1562) );
  NAND3X1 U2170 ( .A(n2323), .B(n2869), .C(n2320), .Y(n2862) );
  NAND4X1 U2171 ( .A(n2855), .B(n2856), .C(n2870), .D(n2871), .Y(n2869) );
  CLKINVX1 U2172 ( .A(a2[8]), .Y(n2868) );
  CLKINVX1 U2173 ( .A(n2874), .Y(n1561) );
  AOI222XL U2174 ( .A0(n2150), .A1(n2875), .B0(n2876), .B1(N1291), .C0(N1291), 
        .C1(n2877), .Y(n2874) );
  CLKINVX1 U2175 ( .A(n2878), .Y(n1560) );
  AOI222XL U2176 ( .A0(n2150), .A1(n2879), .B0(n2876), .B1(max11[1]), .C0(
        N1292), .C1(n2877), .Y(n2878) );
  CLKINVX1 U2177 ( .A(n2880), .Y(n1559) );
  AOI222XL U2178 ( .A0(n2151), .A1(n2881), .B0(n2876), .B1(max11[2]), .C0(
        N1293), .C1(n2877), .Y(n2880) );
  CLKINVX1 U2179 ( .A(n2882), .Y(n1558) );
  AOI222XL U2180 ( .A0(n2150), .A1(n2883), .B0(n2876), .B1(max11[3]), .C0(
        N1294), .C1(n2877), .Y(n2882) );
  CLKINVX1 U2181 ( .A(n2884), .Y(n1557) );
  AOI222XL U2182 ( .A0(n2151), .A1(n2885), .B0(n2876), .B1(max11[4]), .C0(
        N1295), .C1(n2877), .Y(n2884) );
  CLKINVX1 U2183 ( .A(n2886), .Y(n1556) );
  AOI222XL U2184 ( .A0(n2150), .A1(n2887), .B0(n2876), .B1(max11[5]), .C0(
        N1296), .C1(n2877), .Y(n2886) );
  CLKINVX1 U2185 ( .A(n2888), .Y(n1555) );
  AOI222XL U2186 ( .A0(n2151), .A1(n2889), .B0(n2876), .B1(max11[6]), .C0(
        N1297), .C1(n2877), .Y(n2888) );
  CLKINVX1 U2187 ( .A(n2890), .Y(n1554) );
  AOI222XL U2188 ( .A0(n2150), .A1(n2891), .B0(n2876), .B1(max11[7]), .C0(
        N1298), .C1(n2877), .Y(n2890) );
  AO22X1 U2189 ( .A0(a3_8_), .A1(n2152), .B0(n1778), .B1(n2877), .Y(n1553) );
  CLKINVX1 U2190 ( .A(s1), .Y(n2841) );
  CLKINVX1 U2191 ( .A(n2892), .Y(n1552) );
  AOI222XL U2192 ( .A0(n2150), .A1(n2893), .B0(n2894), .B1(N1310), .C0(N1310), 
        .C1(n2895), .Y(n2892) );
  CLKINVX1 U2193 ( .A(n2896), .Y(n1551) );
  AOI222XL U2194 ( .A0(n2151), .A1(n2897), .B0(n2894), .B1(max12[1]), .C0(
        N1311), .C1(n2895), .Y(n2896) );
  CLKINVX1 U2195 ( .A(n2898), .Y(n1550) );
  AOI222XL U2196 ( .A0(n2151), .A1(n2899), .B0(n2894), .B1(max12[2]), .C0(
        N1312), .C1(n2895), .Y(n2898) );
  CLKINVX1 U2197 ( .A(n2900), .Y(n1549) );
  AOI222XL U2198 ( .A0(n2150), .A1(n2901), .B0(n2894), .B1(max12[3]), .C0(
        N1313), .C1(n2895), .Y(n2900) );
  CLKINVX1 U2199 ( .A(n2902), .Y(n1548) );
  AOI222XL U2200 ( .A0(n2150), .A1(n2903), .B0(n2894), .B1(max12[4]), .C0(
        N1314), .C1(n2895), .Y(n2902) );
  CLKINVX1 U2201 ( .A(n2904), .Y(n1547) );
  AOI222XL U2202 ( .A0(n2150), .A1(n2905), .B0(n2894), .B1(max12[5]), .C0(
        N1315), .C1(n2895), .Y(n2904) );
  CLKINVX1 U2203 ( .A(n2906), .Y(n1546) );
  AOI222XL U2204 ( .A0(n2150), .A1(n2907), .B0(n2894), .B1(max12[6]), .C0(
        N1316), .C1(n2895), .Y(n2906) );
  CLKINVX1 U2205 ( .A(n2908), .Y(n1545) );
  AOI222XL U2206 ( .A0(n2150), .A1(n2909), .B0(n2894), .B1(max12[7]), .C0(
        N1317), .C1(n2895), .Y(n2908) );
  AO22X1 U2207 ( .A0(a4_8_), .A1(n2152), .B0(n1779), .B1(n2895), .Y(n1544) );
  CLKINVX1 U2208 ( .A(s2), .Y(n2842) );
  CLKINVX1 U2209 ( .A(n2910), .Y(n1543) );
  AOI222XL U2210 ( .A0(n2150), .A1(n2911), .B0(n2912), .B1(N1329), .C0(N1329), 
        .C1(n2913), .Y(n2910) );
  CLKINVX1 U2211 ( .A(n2914), .Y(n1542) );
  AOI222XL U2212 ( .A0(n2150), .A1(n2915), .B0(n2912), .B1(max21[1]), .C0(
        N1330), .C1(n2913), .Y(n2914) );
  CLKINVX1 U2213 ( .A(n2916), .Y(n1541) );
  AOI222XL U2214 ( .A0(n2150), .A1(n2917), .B0(n2912), .B1(max21[2]), .C0(
        N1331), .C1(n2913), .Y(n2916) );
  CLKINVX1 U2215 ( .A(n2918), .Y(n1540) );
  AOI222XL U2216 ( .A0(n2150), .A1(n2919), .B0(n2912), .B1(max21[3]), .C0(
        N1332), .C1(n2913), .Y(n2918) );
  CLKINVX1 U2217 ( .A(n2920), .Y(n1539) );
  AOI222XL U2218 ( .A0(n2150), .A1(n2921), .B0(n2912), .B1(max21[4]), .C0(
        N1333), .C1(n2913), .Y(n2920) );
  CLKINVX1 U2219 ( .A(n2922), .Y(n1538) );
  AOI222XL U2220 ( .A0(n2150), .A1(n2923), .B0(n2912), .B1(max21[5]), .C0(
        N1334), .C1(n2913), .Y(n2922) );
  CLKINVX1 U2221 ( .A(n2924), .Y(n1537) );
  AOI222XL U2222 ( .A0(n2150), .A1(n2925), .B0(n2912), .B1(max21[6]), .C0(
        N1335), .C1(n2913), .Y(n2924) );
  CLKINVX1 U2223 ( .A(n2926), .Y(n1536) );
  AOI222XL U2224 ( .A0(n2151), .A1(n2927), .B0(n2912), .B1(max21[7]), .C0(
        N1336), .C1(n2913), .Y(n2926) );
  AO22X1 U2225 ( .A0(a5_8_), .A1(n2152), .B0(n1780), .B1(n2913), .Y(n1535) );
  CLKINVX1 U2226 ( .A(s3), .Y(n2843) );
  CLKINVX1 U2227 ( .A(n2928), .Y(n1534) );
  AOI222XL U2228 ( .A0(n2151), .A1(n2929), .B0(n2930), .B1(N1348), .C0(N1348), 
        .C1(n2931), .Y(n2928) );
  CLKINVX1 U2229 ( .A(n2932), .Y(n1533) );
  AOI222XL U2230 ( .A0(n2151), .A1(n2933), .B0(n2930), .B1(max22[1]), .C0(
        N1349), .C1(n2931), .Y(n2932) );
  CLKINVX1 U2231 ( .A(n2934), .Y(n1532) );
  AOI222XL U2232 ( .A0(n2151), .A1(n2935), .B0(n2930), .B1(max22[2]), .C0(
        N1350), .C1(n2931), .Y(n2934) );
  CLKINVX1 U2233 ( .A(n2936), .Y(n1531) );
  AOI222XL U2234 ( .A0(n2151), .A1(n2937), .B0(n2930), .B1(max22[3]), .C0(
        N1351), .C1(n2931), .Y(n2936) );
  CLKINVX1 U2235 ( .A(n2938), .Y(n1530) );
  AOI222XL U2236 ( .A0(n2151), .A1(n2939), .B0(n2930), .B1(max22[4]), .C0(
        N1352), .C1(n2931), .Y(n2938) );
  CLKINVX1 U2237 ( .A(n2940), .Y(n1529) );
  AOI222XL U2238 ( .A0(n2151), .A1(n2941), .B0(n2930), .B1(max22[5]), .C0(
        N1353), .C1(n2931), .Y(n2940) );
  CLKINVX1 U2239 ( .A(n2942), .Y(n1528) );
  AOI222XL U2240 ( .A0(n2151), .A1(n2943), .B0(n2930), .B1(max22[6]), .C0(
        N1354), .C1(n2931), .Y(n2942) );
  CLKINVX1 U2241 ( .A(n2944), .Y(n1527) );
  AOI222XL U2242 ( .A0(n2151), .A1(n2945), .B0(n2930), .B1(max22[7]), .C0(
        N1355), .C1(n2931), .Y(n2944) );
  OAI2BB2XL U2243 ( .B0(n2946), .B1(n2153), .A0N(n1781), .A1N(n2931), .Y(n1526) );
  CLKINVX1 U2244 ( .A(s4), .Y(n2844) );
  CLKINVX1 U2245 ( .A(n2947), .Y(n1525) );
  AOI222XL U2246 ( .A0(n2151), .A1(n2948), .B0(N990), .B1(n2949), .C0(N1402), 
        .C1(n2090), .Y(n2947) );
  CLKINVX1 U2247 ( .A(n2951), .Y(n1524) );
  AOI222XL U2248 ( .A0(n2152), .A1(n2952), .B0(N991), .B1(n2949), .C0(N1403), 
        .C1(n2090), .Y(n2951) );
  CLKINVX1 U2249 ( .A(n2953), .Y(n1523) );
  AOI222XL U2250 ( .A0(n2151), .A1(n2954), .B0(N992), .B1(n2949), .C0(N1404), 
        .C1(n2090), .Y(n2953) );
  CLKINVX1 U2251 ( .A(n2955), .Y(n1522) );
  AOI222XL U2252 ( .A0(n2152), .A1(n2956), .B0(N993), .B1(n2949), .C0(N1405), 
        .C1(n2090), .Y(n2955) );
  CLKINVX1 U2253 ( .A(n2957), .Y(n1521) );
  AOI222XL U2254 ( .A0(n2152), .A1(n2958), .B0(N994), .B1(n2949), .C0(N1406), 
        .C1(n2090), .Y(n2957) );
  CLKINVX1 U2255 ( .A(n2959), .Y(n1520) );
  AOI222XL U2256 ( .A0(n2152), .A1(n2960), .B0(N995), .B1(n2949), .C0(N1407), 
        .C1(n2090), .Y(n2959) );
  CLKINVX1 U2257 ( .A(n2961), .Y(n1519) );
  AOI222XL U2258 ( .A0(n2151), .A1(n2962), .B0(N996), .B1(n2949), .C0(N1408), 
        .C1(n2090), .Y(n2961) );
  CLKINVX1 U2259 ( .A(n2963), .Y(n1518) );
  AOI222XL U2260 ( .A0(n2151), .A1(n2964), .B0(N997), .B1(n2949), .C0(N1409), 
        .C1(n2090), .Y(n2963) );
  OAI2BB2XL U2261 ( .B0(n1697), .B1(n745), .A0N(N1410), .A1N(n2090), .Y(n1517)
         );
  XOR3X1 U2262 ( .A(n2966), .B(n2967), .C(n2968), .Y(n2965) );
  OAI22XL U2263 ( .A0(n2817), .A1(n2203), .B0(n2969), .B1(n2970), .Y(n2968) );
  OAI32X1 U2264 ( .A0(n2972), .A1(n2332), .A2(n2345), .B0(n2973), .B1(n2331), 
        .Y(n1516) );
  CLKINVX1 U2265 ( .A(a1[0]), .Y(n2331) );
  CLKINVX1 U2266 ( .A(n2974), .Y(n2973) );
  AOI211X1 U2267 ( .A0(n2975), .A1(a1[0]), .B0(n2976), .C0(n2977), .Y(n2332)
         );
  CLKMX2X2 U2268 ( .A(n2978), .B(n2979), .S0(node[0]), .Y(n2977) );
  OAI21XL U2269 ( .A0(n2853), .A1(n2326), .B0(n2855), .Y(n2979) );
  NAND2BX1 U2270 ( .AN(n2980), .B(n2981), .Y(n2855) );
  CLKINVX1 U2271 ( .A(n2982), .Y(n2326) );
  OAI21XL U2272 ( .A0(n2983), .A1(n2872), .B0(n2859), .Y(n2978) );
  CLKINVX1 U2273 ( .A(n2984), .Y(n1515) );
  OAI21XL U2274 ( .A0(n2333), .A1(n2177), .B0(n2986), .Y(n2974) );
  NAND4X1 U2275 ( .A(n2987), .B(n2856), .C(n2988), .D(n2989), .Y(n2344) );
  AOI221XL U2276 ( .A0(n2982), .A1(n2990), .B0(a1[1]), .B1(n2975), .C0(n2976), 
        .Y(n2989) );
  OR2X1 U2277 ( .A(n2853), .B(n2980), .Y(n2988) );
  NAND2X1 U2278 ( .A(node[1]), .B(n2872), .Y(n2853) );
  OAI2BB1X1 U2279 ( .A0N(n2859), .A1N(n2983), .B0(node[0]), .Y(n2987) );
  NAND3X1 U2280 ( .A(node[4]), .B(node[3]), .C(n2981), .Y(n2859) );
  OAI21XL U2281 ( .A0(n786), .A1(n2991), .B0(n2992), .Y(n1514) );
  OAI21XL U2282 ( .A0(n785), .A1(n2991), .B0(n2992), .Y(n1513) );
  OAI21XL U2283 ( .A0(n784), .A1(n2991), .B0(n2992), .Y(n1512) );
  OAI21XL U2284 ( .A0(n783), .A1(n2991), .B0(n2992), .Y(n1511) );
  OAI21XL U2285 ( .A0(n782), .A1(n2991), .B0(n2992), .Y(n1510) );
  OAI21XL U2286 ( .A0(n781), .A1(n2991), .B0(n2992), .Y(n1509) );
  OAI21XL U2287 ( .A0(n780), .A1(n2991), .B0(n2992), .Y(n1508) );
  NAND2X1 U2288 ( .A(n2993), .B(n2985), .Y(n2992) );
  CLKINVX1 U2289 ( .A(n2972), .Y(n2985) );
  OAI21XL U2290 ( .A0(n2996), .A1(n2997), .B0(n2172), .Y(n2995) );
  OA21XL U2291 ( .A0(n786), .A1(n2873), .B0(n3002), .Y(n3001) );
  AOI211X1 U2292 ( .A0(a2[2]), .A1(n2092), .B0(n3004), .C0(n3005), .Y(n2998)
         );
  OAI22XL U2293 ( .A0(n777), .A1(n2337), .B0(n751), .B1(n2338), .Y(n3005) );
  OAI222XL U2294 ( .A0(n740), .A1(n2339), .B0(n759), .B1(n2340), .C0(n768), 
        .C1(n2341), .Y(n3004) );
  OA21XL U2295 ( .A0(n785), .A1(n2873), .B0(n3002), .Y(n3008) );
  AOI211X1 U2296 ( .A0(a2[3]), .A1(n2092), .B0(n3009), .C0(n3010), .Y(n3006)
         );
  OAI22XL U2297 ( .A0(n776), .A1(n2337), .B0(n750), .B1(n2338), .Y(n3010) );
  OAI222XL U2298 ( .A0(n739), .A1(n2339), .B0(n758), .B1(n2340), .C0(n767), 
        .C1(n2341), .Y(n3009) );
  OA21XL U2299 ( .A0(n784), .A1(n2873), .B0(n3002), .Y(n3013) );
  AOI211X1 U2300 ( .A0(a2[4]), .A1(n2092), .B0(n3014), .C0(n3015), .Y(n3011)
         );
  OAI22XL U2301 ( .A0(n775), .A1(n2337), .B0(n749), .B1(n2338), .Y(n3015) );
  OAI222XL U2302 ( .A0(n738), .A1(n2339), .B0(n757), .B1(n2340), .C0(n766), 
        .C1(n2341), .Y(n3014) );
  OA21XL U2303 ( .A0(n783), .A1(n2873), .B0(n3002), .Y(n3018) );
  AOI211X1 U2304 ( .A0(a2[5]), .A1(n2092), .B0(n3019), .C0(n3020), .Y(n3016)
         );
  OAI22XL U2305 ( .A0(n774), .A1(n2337), .B0(n748), .B1(n2338), .Y(n3020) );
  OAI222XL U2306 ( .A0(n737), .A1(n2339), .B0(n756), .B1(n2340), .C0(n765), 
        .C1(n2341), .Y(n3019) );
  OA21XL U2307 ( .A0(n782), .A1(n2873), .B0(n3002), .Y(n3023) );
  AOI211X1 U2308 ( .A0(a2[6]), .A1(n2092), .B0(n3024), .C0(n3025), .Y(n3021)
         );
  OAI22XL U2309 ( .A0(n773), .A1(n2337), .B0(n747), .B1(n2338), .Y(n3025) );
  OAI222XL U2310 ( .A0(n736), .A1(n2339), .B0(n755), .B1(n2340), .C0(n764), 
        .C1(n2341), .Y(n3024) );
  OAI211X1 U2311 ( .A0(n3026), .A1(n2999), .B0(n3027), .C0(n3028), .Y(n1502)
         );
  OA21XL U2312 ( .A0(n781), .A1(n2873), .B0(n3002), .Y(n3028) );
  AOI211X1 U2313 ( .A0(a2[7]), .A1(n2092), .B0(n3029), .C0(n3030), .Y(n3026)
         );
  OAI22XL U2314 ( .A0(n772), .A1(n2337), .B0(n746), .B1(n2338), .Y(n3030) );
  OAI222XL U2315 ( .A0(n735), .A1(n2339), .B0(n754), .B1(n2340), .C0(n763), 
        .C1(n2341), .Y(n3029) );
  OA21XL U2316 ( .A0(n780), .A1(n2873), .B0(n3002), .Y(n3035) );
  NAND2X1 U2317 ( .A(n2993), .B(n2323), .Y(n3002) );
  CLKINVX1 U2318 ( .A(n3036), .Y(n2993) );
  OAI31XL U2319 ( .A0(n3037), .A1(n3038), .A2(n2976), .B0(n2333), .Y(n3036) );
  CLKMX2X2 U2320 ( .A(n3039), .B(n3040), .S0(node[0]), .Y(n2976) );
  OAI2BB1X1 U2321 ( .A0N(n2981), .A1N(n2982), .B0(n2856), .Y(n3040) );
  OAI221XL U2322 ( .A0(n2980), .A1(n2324), .B0(n2990), .B1(n2858), .C0(n2860), 
        .Y(n3039) );
  NAND3X1 U2323 ( .A(node[2]), .B(node[1]), .C(n2982), .Y(n2860) );
  CLKINVX1 U2324 ( .A(node[2]), .Y(n2872) );
  OA21XL U2325 ( .A0(n2851), .A1(n2981), .B0(n2982), .Y(n3038) );
  NOR2X1 U2326 ( .A(n2325), .B(node[3]), .Y(n2982) );
  NOR2X1 U2327 ( .A(n2857), .B(n2324), .Y(n2851) );
  NAND2X1 U2328 ( .A(node[2]), .B(n2990), .Y(n2324) );
  OAI31XL U2329 ( .A0(n2857), .A1(node[2]), .A2(n2983), .B0(n2856), .Y(n3037)
         );
  NAND4X1 U2330 ( .A(node[2]), .B(node[1]), .C(n2850), .D(n2325), .Y(n2856) );
  AOI2BB1X1 U2331 ( .A0N(n2990), .A1N(n2980), .B0(n2852), .Y(n2983) );
  CLKINVX1 U2332 ( .A(n2870), .Y(n2852) );
  NAND2X1 U2333 ( .A(node[3]), .B(n2325), .Y(n2980) );
  CLKINVX1 U2334 ( .A(node[0]), .Y(n2857) );
  NOR2X1 U2335 ( .A(n2345), .B(n2975), .Y(n2994) );
  OAI33X1 U2336 ( .A0(n2870), .A1(node[2]), .A2(node[0]), .B0(n2325), .B1(
        n2981), .B2(n2850), .Y(n2975) );
  NOR2X1 U2337 ( .A(node[1]), .B(node[2]), .Y(n2981) );
  CLKINVX1 U2338 ( .A(node[1]), .Y(n2990) );
  CLKINVX1 U2339 ( .A(node[3]), .Y(n2850) );
  NAND2X1 U2340 ( .A(n3041), .B(n8330), .Y(n2999) );
  NOR4BX1 U2341 ( .AN(n3044), .B(N1077), .C(N1076), .D(n2328), .Y(n3043) );
  NOR3X1 U2342 ( .A(N1078), .B(N1080), .C(N1079), .Y(n3044) );
  OR4X1 U2343 ( .A(n3045), .B(n3031), .C(n2092), .D(n3032), .Y(n3042) );
  NAND3X1 U2344 ( .A(n2338), .B(n2337), .C(n2341), .Y(n3045) );
  AOI211X1 U2345 ( .A0(a2[8]), .A1(n2092), .B0(n3046), .C0(n3047), .Y(n3033)
         );
  OAI22XL U2346 ( .A0(n2337), .A1(n2946), .B0(n745), .B1(n2338), .Y(n3047) );
  CLKINVX1 U2347 ( .A(a6_8_), .Y(n2946) );
  CLKINVX1 U2348 ( .A(n3049), .Y(n3046) );
  AOI222XL U2349 ( .A0(n3032), .A1(a3_8_), .B0(n3031), .B1(a4_8_), .C0(n3050), 
        .C1(a5_8_), .Y(n3049) );
  CLKINVX1 U2350 ( .A(n2341), .Y(n3050) );
  NOR3X1 U2351 ( .A(N1075), .B(outmode[0]), .C(n3048), .Y(n3031) );
  NOR3X1 U2352 ( .A(N1073), .B(N1075), .C(n3048), .Y(n3032) );
  CLKINVX1 U2353 ( .A(N1074), .Y(n3048) );
  NOR3X1 U2354 ( .A(N1075), .B(outmode[0]), .C(N1074), .Y(n2334) );
  NOR2X1 U2355 ( .A(n3051), .B(n2804), .Y(n2350) );
  CLKINVX1 U2356 ( .A(n2783), .Y(n2367) );
  NOR2X1 U2357 ( .A(n2803), .B(N1001), .Y(n2783) );
  NAND2X1 U2358 ( .A(n3059), .B(N1001), .Y(n2793) );
  NAND2X1 U2359 ( .A(n3059), .B(mode[0]), .Y(n2794) );
  NOR2X1 U2360 ( .A(mode[2]), .B(n390), .Y(n3059) );
  NAND2X1 U2361 ( .A(n3060), .B(N1001), .Y(n2795) );
  NAND2X1 U2362 ( .A(n3060), .B(mode[0]), .Y(n2791) );
  NOR2X1 U2363 ( .A(mode[1]), .B(n388), .Y(n3060) );
  NAND2X1 U2364 ( .A(n3061), .B(N1001), .Y(n2790) );
  NOR2X1 U2365 ( .A(n388), .B(n390), .Y(n3061) );
  NAND4X1 U2366 ( .A(n2792), .B(n2365), .C(n2351), .D(n2801), .Y(n3063) );
  NAND2X1 U2367 ( .A(n390), .B(n388), .Y(n2803) );
  NAND2X1 U2368 ( .A(in_valid), .B(n2170), .Y(n2348) );
  NOR3X1 U2369 ( .A(n383), .B(n386), .C(mode[4]), .Y(n2792) );
  CLKINVX1 U2370 ( .A(n2840), .Y(N937) );
  CLKINVX1 U2371 ( .A(n2838), .Y(N935) );
  CLKINVX1 U2372 ( .A(n2837), .Y(N934) );
  CLKINVX1 U2373 ( .A(n2836), .Y(N933) );
  CLKINVX1 U2374 ( .A(n2835), .Y(N932) );
  CLKINVX1 U2375 ( .A(n2834), .Y(N931) );
  MXI2X1 U2376 ( .A(N923), .B(N915), .S0(n2088), .Y(n2834) );
  CLKINVX1 U2377 ( .A(n2832), .Y(N910) );
  MXI2X1 U2378 ( .A(N901), .B(N893), .S0(N885), .Y(n2831) );
  CLKINVX1 U2379 ( .A(n2830), .Y(N908) );
  MXI2X1 U2380 ( .A(N900), .B(N892), .S0(N885), .Y(n2830) );
  CLKINVX1 U2381 ( .A(n2829), .Y(N907) );
  MXI2X1 U2382 ( .A(N899), .B(N891), .S0(N885), .Y(n2829) );
  CLKINVX1 U2383 ( .A(n2828), .Y(N906) );
  MXI2X1 U2384 ( .A(N898), .B(N890), .S0(N885), .Y(n2828) );
  CLKINVX1 U2385 ( .A(n2827), .Y(N905) );
  MXI2X1 U2386 ( .A(N897), .B(N889), .S0(N885), .Y(n2827) );
  MXI2X1 U2387 ( .A(N875), .B(N867), .S0(N858), .Y(n2824) );
  MXI2X1 U2388 ( .A(N874), .B(N866), .S0(N858), .Y(n2823) );
  MXI2X1 U2389 ( .A(N873), .B(N865), .S0(N858), .Y(n2822) );
  MXI2X1 U2390 ( .A(N872), .B(N864), .S0(N858), .Y(n2821) );
  MXI2X1 U2391 ( .A(N871), .B(N863), .S0(N858), .Y(n2820) );
  MXI2X1 U2392 ( .A(N870), .B(N862), .S0(N858), .Y(n2819) );
  CLKINVX1 U2393 ( .A(n2818), .Y(N877) );
  MXI2X1 U2394 ( .A(N869), .B(N861), .S0(N858), .Y(n2818) );
  MXI2X1 U2395 ( .A(N848), .B(N840), .S0(n1777), .Y(n2815) );
  MXI2X1 U2396 ( .A(N847), .B(N839), .S0(n1777), .Y(n2814) );
  MXI2X1 U2397 ( .A(N846), .B(N838), .S0(n1777), .Y(n2813) );
  MXI2X1 U2398 ( .A(N843), .B(N835), .S0(n1777), .Y(n2810) );
  CLKINVX1 U2399 ( .A(n2809), .Y(N850) );
  OAI2BB1X1 U2400 ( .A0N(n3064), .A1N(n2173), .B0(n3065), .Y(N183) );
  OAI21XL U2401 ( .A0(n3056), .A1(n3066), .B0(n3041), .Y(n3065) );
  NAND2X1 U2402 ( .A(n2316), .B(n3068), .Y(n3064) );
  OAI21XL U2403 ( .A0(mode[2]), .A1(n2804), .B0(n2785), .Y(n3068) );
  CLKINVX1 U2404 ( .A(n2784), .Y(n2804) );
  NOR2X1 U2405 ( .A(n2352), .B(n2177), .Y(n3041) );
  CLKINVX1 U2406 ( .A(n2094), .Y(n2352) );
  NOR3X1 U2407 ( .A(n2179), .B(n3066), .C(n3056), .Y(n3067) );
  NOR2X1 U2408 ( .A(n3051), .B(mode[5]), .Y(n3056) );
  CLKINVX1 U2409 ( .A(n3069), .Y(n3066) );
  OAI211X1 U2410 ( .A0(n386), .A1(n388), .B0(n3070), .C0(n3071), .Y(n3069) );
  NOR2X1 U2411 ( .A(mode[4]), .B(n3051), .Y(n3071) );
  CLKINVX1 U2412 ( .A(n2801), .Y(n3051) );
  NOR2X1 U2413 ( .A(n2785), .B(mode[7]), .Y(n2801) );
  OAI21XL U2414 ( .A0(mode[1]), .A1(mode[0]), .B0(mode[3]), .Y(n3070) );
endmodule

